##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Tue Apr 20 14:00:48 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_single2
  CLASS BLOCK ;
  SIZE 230.4600 BY 30.2600 ;
  FOREIGN S_term_single2 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.0050 29.9300 19.1750 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.6250 29.9300 17.7950 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.2450 29.9300 16.4150 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.3250 29.9300 15.4950 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 29.5850 29.9300 29.7550 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 28.2050 29.9300 28.3750 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 26.8250 29.9300 26.9950 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.9050 29.9300 26.0750 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.5250 29.9300 24.6950 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.1450 29.9300 23.3150 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.7650 29.9300 21.9350 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 20.3850 29.9300 20.5550 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 40.1650 29.9300 40.3350 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 38.7850 29.9300 38.9550 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 37.8650 29.9300 38.0350 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 36.4850 29.9300 36.6550 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 35.1050 29.9300 35.2750 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 33.7250 29.9300 33.8950 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 32.3450 29.9300 32.5150 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 30.9650 29.9300 31.1350 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 61.7850 29.9300 61.9550 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 60.4050 29.9300 60.5750 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 59.0250 29.9300 59.1950 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 57.6450 29.9300 57.8150 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 56.2650 29.9300 56.4350 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 54.8850 29.9300 55.0550 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 53.5050 29.9300 53.6750 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 52.1250 29.9300 52.2950 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 50.7450 29.9300 50.9150 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 49.8250 29.9300 49.9950 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 48.4450 29.9300 48.6150 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 47.0650 29.9300 47.2350 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 45.6850 29.9300 45.8550 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 44.3050 29.9300 44.4750 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 42.9250 29.9300 43.0950 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 41.5450 29.9300 41.7150 30.2600 ;
    END
  END N4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 66.8450 29.9300 67.0150 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 65.4650 29.9300 65.6350 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 64.0850 29.9300 64.2550 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 62.7050 29.9300 62.8750 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 88.0050 29.9300 88.1750 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 86.6250 29.9300 86.7950 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 85.7050 29.9300 85.8750 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 84.3250 29.9300 84.4950 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 82.9450 29.9300 83.1150 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 81.5650 29.9300 81.7350 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 80.1850 29.9300 80.3550 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 78.8050 29.9300 78.9750 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 77.4250 29.9300 77.5950 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 76.0450 29.9300 76.2150 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 74.6650 29.9300 74.8350 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 73.7450 29.9300 73.9150 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 72.3650 29.9300 72.5350 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 70.9850 29.9300 71.1550 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 69.6050 29.9300 69.7750 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 68.2250 29.9300 68.3950 30.2600 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 109.6250 29.9300 109.7950 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 108.2450 29.9300 108.4150 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 106.8650 29.9300 107.0350 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 105.4850 29.9300 105.6550 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 104.1050 29.9300 104.2750 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 102.7250 29.9300 102.8950 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 101.3450 29.9300 101.5150 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 99.9650 29.9300 100.1350 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 98.5850 29.9300 98.7550 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 97.6650 29.9300 97.8350 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 96.2850 29.9300 96.4550 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 94.9050 29.9300 95.0750 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 93.5250 29.9300 93.6950 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 92.1450 29.9300 92.3150 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 90.7650 29.9300 90.9350 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 89.3850 29.9300 89.5550 30.2600 ;
    END
  END S4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 26.6800 0.8000 26.9800 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 24.8500 0.8000 25.1500 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 23.0200 0.8000 23.3200 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 21.8000 0.8000 22.1000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 19.9700 0.8000 20.2700 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 18.7500 0.8000 19.0500 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 16.9200 0.8000 17.2200 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 15.0900 0.8000 15.3900 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 13.8700 0.8000 14.1700 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 12.0400 0.8000 12.3400 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 10.8200 0.8000 11.1200 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 8.9900 0.8000 9.2900 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 7.1600 0.8000 7.4600 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 5.9400 0.8000 6.2400 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 4.1100 0.8000 4.4100 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2.8900 0.8000 3.1900 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 27.6400 0.5950 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.9400 0.5950 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 24.2400 0.5950 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.5400 0.5950 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 20.8400 0.5950 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 19.1400 0.5950 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 17.4400 0.5950 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 15.7400 0.5950 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 14.0400 0.5950 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 12.3400 0.5950 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 10.6400 0.5950 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 8.9400 0.5950 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 7.2400 0.5950 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 5.5400 0.5950 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3.8400 0.5950 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2.1400 0.5950 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 26.6800 230.4600 26.9800 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 24.8500 230.4600 25.1500 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 23.0200 230.4600 23.3200 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 21.8000 230.4600 22.1000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 19.9700 230.4600 20.2700 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 18.7500 230.4600 19.0500 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 16.9200 230.4600 17.2200 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 15.0900 230.4600 15.3900 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 13.8700 230.4600 14.1700 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 12.0400 230.4600 12.3400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 10.8200 230.4600 11.1200 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 8.9900 230.4600 9.2900 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 7.1600 230.4600 7.4600 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 5.9400 230.4600 6.2400 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 4.1100 230.4600 4.4100 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.6600 2.8900 230.4600 3.1900 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 27.6400 230.4600 27.7800 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 25.9400 230.4600 26.0800 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 24.2400 230.4600 24.3800 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 22.5400 230.4600 22.6800 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 20.8400 230.4600 20.9800 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 19.1400 230.4600 19.2800 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 17.4400 230.4600 17.5800 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 15.7400 230.4600 15.8800 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 14.0400 230.4600 14.1800 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 12.3400 230.4600 12.4800 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 10.6400 230.4600 10.7800 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 8.9400 230.4600 9.0800 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 7.2400 230.4600 7.3800 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 5.5400 230.4600 5.6800 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 3.8400 230.4600 3.9800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 229.8650 2.1400 230.4600 2.2800 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.0600 0.0000 214.2000 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.4600 0.0000 209.6000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.4000 0.0000 204.5400 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.3400 0.0000 199.4800 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.2800 0.0000 194.4200 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.6800 0.0000 189.8200 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.6200 0.0000 184.7600 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.5600 0.0000 179.7000 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.5000 0.0000 174.6400 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.4400 0.0000 169.5800 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.8400 0.0000 164.9800 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.7800 0.0000 159.9200 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.7200 0.0000 154.8600 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.6600 0.0000 149.8000 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.6000 0.0000 144.7400 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.0000 0.0000 140.1400 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.9400 0.0000 135.0800 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.8800 0.0000 130.0200 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.8200 0.0000 124.9600 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.2200 0.0000 120.3600 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.0600 29.7750 214.2000 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.4600 29.7750 209.6000 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.4000 29.7750 204.5400 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.3400 29.7750 199.4800 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.2800 29.7750 194.4200 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.6800 29.7750 189.8200 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.6200 29.7750 184.7600 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.5600 29.7750 179.7000 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.5000 29.7750 174.6400 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.4400 29.7750 169.5800 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.8400 29.7750 164.9800 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.7800 29.7750 159.9200 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.7200 29.7750 154.8600 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.6600 29.7750 149.8000 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.6000 29.7750 144.7400 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.0000 29.7750 140.1400 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.9400 29.7750 135.0800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.8800 29.7750 130.0200 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.8200 29.7750 124.9600 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.2200 29.7750 120.3600 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 222.9000 4.0700 224.9000 25.0000 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
      LAYER met3 ;
        RECT 5.5600 4.0700 224.9000 6.0700 ;
        RECT 5.5600 23.0000 224.9000 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 225.9000 1.0700 227.9000 28.0000 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
      LAYER met3 ;
        RECT 2.5600 1.0700 227.9000 3.0700 ;
        RECT 2.5600 26.0000 227.9000 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 109.9650 29.7600 230.4600 30.2600 ;
      RECT 108.5850 29.7600 109.4550 30.2600 ;
      RECT 107.2050 29.7600 108.0750 30.2600 ;
      RECT 105.8250 29.7600 106.6950 30.2600 ;
      RECT 104.4450 29.7600 105.3150 30.2600 ;
      RECT 103.0650 29.7600 103.9350 30.2600 ;
      RECT 101.6850 29.7600 102.5550 30.2600 ;
      RECT 100.3050 29.7600 101.1750 30.2600 ;
      RECT 98.9250 29.7600 99.7950 30.2600 ;
      RECT 98.0050 29.7600 98.4150 30.2600 ;
      RECT 96.6250 29.7600 97.4950 30.2600 ;
      RECT 95.2450 29.7600 96.1150 30.2600 ;
      RECT 93.8650 29.7600 94.7350 30.2600 ;
      RECT 92.4850 29.7600 93.3550 30.2600 ;
      RECT 91.1050 29.7600 91.9750 30.2600 ;
      RECT 89.7250 29.7600 90.5950 30.2600 ;
      RECT 88.3450 29.7600 89.2150 30.2600 ;
      RECT 86.9650 29.7600 87.8350 30.2600 ;
      RECT 86.0450 29.7600 86.4550 30.2600 ;
      RECT 84.6650 29.7600 85.5350 30.2600 ;
      RECT 83.2850 29.7600 84.1550 30.2600 ;
      RECT 81.9050 29.7600 82.7750 30.2600 ;
      RECT 80.5250 29.7600 81.3950 30.2600 ;
      RECT 79.1450 29.7600 80.0150 30.2600 ;
      RECT 77.7650 29.7600 78.6350 30.2600 ;
      RECT 76.3850 29.7600 77.2550 30.2600 ;
      RECT 75.0050 29.7600 75.8750 30.2600 ;
      RECT 74.0850 29.7600 74.4950 30.2600 ;
      RECT 72.7050 29.7600 73.5750 30.2600 ;
      RECT 71.3250 29.7600 72.1950 30.2600 ;
      RECT 69.9450 29.7600 70.8150 30.2600 ;
      RECT 68.5650 29.7600 69.4350 30.2600 ;
      RECT 67.1850 29.7600 68.0550 30.2600 ;
      RECT 65.8050 29.7600 66.6750 30.2600 ;
      RECT 64.4250 29.7600 65.2950 30.2600 ;
      RECT 63.0450 29.7600 63.9150 30.2600 ;
      RECT 62.1250 29.7600 62.5350 30.2600 ;
      RECT 60.7450 29.7600 61.6150 30.2600 ;
      RECT 59.3650 29.7600 60.2350 30.2600 ;
      RECT 57.9850 29.7600 58.8550 30.2600 ;
      RECT 56.6050 29.7600 57.4750 30.2600 ;
      RECT 55.2250 29.7600 56.0950 30.2600 ;
      RECT 53.8450 29.7600 54.7150 30.2600 ;
      RECT 52.4650 29.7600 53.3350 30.2600 ;
      RECT 51.0850 29.7600 51.9550 30.2600 ;
      RECT 50.1650 29.7600 50.5750 30.2600 ;
      RECT 48.7850 29.7600 49.6550 30.2600 ;
      RECT 47.4050 29.7600 48.2750 30.2600 ;
      RECT 46.0250 29.7600 46.8950 30.2600 ;
      RECT 44.6450 29.7600 45.5150 30.2600 ;
      RECT 43.2650 29.7600 44.1350 30.2600 ;
      RECT 41.8850 29.7600 42.7550 30.2600 ;
      RECT 40.5050 29.7600 41.3750 30.2600 ;
      RECT 39.1250 29.7600 39.9950 30.2600 ;
      RECT 38.2050 29.7600 38.6150 30.2600 ;
      RECT 36.8250 29.7600 37.6950 30.2600 ;
      RECT 35.4450 29.7600 36.3150 30.2600 ;
      RECT 34.0650 29.7600 34.9350 30.2600 ;
      RECT 32.6850 29.7600 33.5550 30.2600 ;
      RECT 31.3050 29.7600 32.1750 30.2600 ;
      RECT 29.9250 29.7600 30.7950 30.2600 ;
      RECT 28.5450 29.7600 29.4150 30.2600 ;
      RECT 27.1650 29.7600 28.0350 30.2600 ;
      RECT 26.2450 29.7600 26.6550 30.2600 ;
      RECT 24.8650 29.7600 25.7350 30.2600 ;
      RECT 23.4850 29.7600 24.3550 30.2600 ;
      RECT 22.1050 29.7600 22.9750 30.2600 ;
      RECT 20.7250 29.7600 21.5950 30.2600 ;
      RECT 19.3450 29.7600 20.2150 30.2600 ;
      RECT 17.9650 29.7600 18.8350 30.2600 ;
      RECT 16.5850 29.7600 17.4550 30.2600 ;
      RECT 15.6650 29.7600 16.0750 30.2600 ;
      RECT 0.0000 29.7600 15.1550 30.2600 ;
      RECT 0.0000 0.0000 230.4600 29.7600 ;
    LAYER met1 ;
      RECT 0.0000 27.9200 230.4600 30.2600 ;
      RECT 0.7350 27.5000 229.7250 27.9200 ;
      RECT 0.0000 26.2200 230.4600 27.5000 ;
      RECT 0.7350 25.8000 229.7250 26.2200 ;
      RECT 0.0000 24.5200 230.4600 25.8000 ;
      RECT 0.7350 24.1000 229.7250 24.5200 ;
      RECT 0.0000 22.8200 230.4600 24.1000 ;
      RECT 0.7350 22.4000 229.7250 22.8200 ;
      RECT 0.0000 21.1200 230.4600 22.4000 ;
      RECT 0.7350 20.7000 229.7250 21.1200 ;
      RECT 0.0000 19.4200 230.4600 20.7000 ;
      RECT 0.7350 19.0000 229.7250 19.4200 ;
      RECT 0.0000 17.7200 230.4600 19.0000 ;
      RECT 0.7350 17.3000 229.7250 17.7200 ;
      RECT 0.0000 16.0200 230.4600 17.3000 ;
      RECT 0.7350 15.6000 229.7250 16.0200 ;
      RECT 0.0000 14.3200 230.4600 15.6000 ;
      RECT 0.7350 13.9000 229.7250 14.3200 ;
      RECT 0.0000 12.6200 230.4600 13.9000 ;
      RECT 0.7350 12.2000 229.7250 12.6200 ;
      RECT 0.0000 10.9200 230.4600 12.2000 ;
      RECT 0.7350 10.5000 229.7250 10.9200 ;
      RECT 0.0000 9.2200 230.4600 10.5000 ;
      RECT 0.7350 8.8000 229.7250 9.2200 ;
      RECT 0.0000 7.5200 230.4600 8.8000 ;
      RECT 0.7350 7.1000 229.7250 7.5200 ;
      RECT 0.0000 5.8200 230.4600 7.1000 ;
      RECT 0.7350 5.4000 229.7250 5.8200 ;
      RECT 0.0000 4.1200 230.4600 5.4000 ;
      RECT 0.7350 3.7000 229.7250 4.1200 ;
      RECT 0.0000 2.4200 230.4600 3.7000 ;
      RECT 0.7350 2.0000 229.7250 2.4200 ;
      RECT 0.0000 0.0000 230.4600 2.0000 ;
    LAYER met2 ;
      RECT 214.3400 29.6350 230.4600 30.2600 ;
      RECT 209.7400 29.6350 213.9200 30.2600 ;
      RECT 204.6800 29.6350 209.3200 30.2600 ;
      RECT 199.6200 29.6350 204.2600 30.2600 ;
      RECT 194.5600 29.6350 199.2000 30.2600 ;
      RECT 189.9600 29.6350 194.1400 30.2600 ;
      RECT 184.9000 29.6350 189.5400 30.2600 ;
      RECT 179.8400 29.6350 184.4800 30.2600 ;
      RECT 174.7800 29.6350 179.4200 30.2600 ;
      RECT 169.7200 29.6350 174.3600 30.2600 ;
      RECT 165.1200 29.6350 169.3000 30.2600 ;
      RECT 160.0600 29.6350 164.7000 30.2600 ;
      RECT 155.0000 29.6350 159.6400 30.2600 ;
      RECT 149.9400 29.6350 154.5800 30.2600 ;
      RECT 144.8800 29.6350 149.5200 30.2600 ;
      RECT 140.2800 29.6350 144.4600 30.2600 ;
      RECT 135.2200 29.6350 139.8600 30.2600 ;
      RECT 130.1600 29.6350 134.8000 30.2600 ;
      RECT 125.1000 29.6350 129.7400 30.2600 ;
      RECT 120.5000 29.6350 124.6800 30.2600 ;
      RECT 0.0000 29.6350 120.0800 30.2600 ;
      RECT 0.0000 28.1400 230.4600 29.6350 ;
      RECT 4.7000 25.1400 225.7600 28.1400 ;
      RECT 225.0400 3.9300 225.7600 25.1400 ;
      RECT 7.7000 3.9300 222.7600 25.1400 ;
      RECT 4.7000 3.9300 5.4200 25.1400 ;
      RECT 228.0400 0.9300 230.4600 28.1400 ;
      RECT 4.7000 0.9300 225.7600 3.9300 ;
      RECT 0.0000 0.9300 2.4200 28.1400 ;
      RECT 0.0000 0.6250 230.4600 0.9300 ;
      RECT 214.3400 0.0000 230.4600 0.6250 ;
      RECT 209.7400 0.0000 213.9200 0.6250 ;
      RECT 204.6800 0.0000 209.3200 0.6250 ;
      RECT 199.6200 0.0000 204.2600 0.6250 ;
      RECT 194.5600 0.0000 199.2000 0.6250 ;
      RECT 189.9600 0.0000 194.1400 0.6250 ;
      RECT 184.9000 0.0000 189.5400 0.6250 ;
      RECT 179.8400 0.0000 184.4800 0.6250 ;
      RECT 174.7800 0.0000 179.4200 0.6250 ;
      RECT 169.7200 0.0000 174.3600 0.6250 ;
      RECT 165.1200 0.0000 169.3000 0.6250 ;
      RECT 160.0600 0.0000 164.7000 0.6250 ;
      RECT 155.0000 0.0000 159.6400 0.6250 ;
      RECT 149.9400 0.0000 154.5800 0.6250 ;
      RECT 144.8800 0.0000 149.5200 0.6250 ;
      RECT 140.2800 0.0000 144.4600 0.6250 ;
      RECT 135.2200 0.0000 139.8600 0.6250 ;
      RECT 130.1600 0.0000 134.8000 0.6250 ;
      RECT 125.1000 0.0000 129.7400 0.6250 ;
      RECT 120.5000 0.0000 124.6800 0.6250 ;
      RECT 0.0000 0.0000 120.0800 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 230.4600 30.2600 ;
      RECT 228.2000 27.2800 230.4600 28.3000 ;
      RECT 0.0000 27.2800 2.2600 28.3000 ;
      RECT 228.2000 26.3800 229.3600 27.2800 ;
      RECT 1.1000 26.3800 2.2600 27.2800 ;
      RECT 228.2000 25.7000 230.4600 26.3800 ;
      RECT 0.0000 25.7000 2.2600 26.3800 ;
      RECT 0.0000 25.4500 230.4600 25.7000 ;
      RECT 1.1000 25.3000 229.3600 25.4500 ;
      RECT 225.2000 24.5500 229.3600 25.3000 ;
      RECT 1.1000 24.5500 5.2600 25.3000 ;
      RECT 225.2000 23.6200 230.4600 24.5500 ;
      RECT 0.0000 23.6200 5.2600 24.5500 ;
      RECT 225.2000 22.7200 229.3600 23.6200 ;
      RECT 1.1000 22.7200 5.2600 23.6200 ;
      RECT 225.2000 22.7000 230.4600 22.7200 ;
      RECT 0.0000 22.7000 5.2600 22.7200 ;
      RECT 0.0000 22.4000 230.4600 22.7000 ;
      RECT 1.1000 21.5000 229.3600 22.4000 ;
      RECT 0.0000 20.5700 230.4600 21.5000 ;
      RECT 1.1000 19.6700 229.3600 20.5700 ;
      RECT 0.0000 19.3500 230.4600 19.6700 ;
      RECT 1.1000 18.4500 229.3600 19.3500 ;
      RECT 0.0000 17.5200 230.4600 18.4500 ;
      RECT 1.1000 16.6200 229.3600 17.5200 ;
      RECT 0.0000 15.6900 230.4600 16.6200 ;
      RECT 1.1000 14.7900 229.3600 15.6900 ;
      RECT 0.0000 14.4700 230.4600 14.7900 ;
      RECT 1.1000 13.5700 229.3600 14.4700 ;
      RECT 0.0000 12.6400 230.4600 13.5700 ;
      RECT 1.1000 11.7400 229.3600 12.6400 ;
      RECT 0.0000 11.4200 230.4600 11.7400 ;
      RECT 1.1000 10.5200 229.3600 11.4200 ;
      RECT 0.0000 9.5900 230.4600 10.5200 ;
      RECT 1.1000 8.6900 229.3600 9.5900 ;
      RECT 0.0000 7.7600 230.4600 8.6900 ;
      RECT 1.1000 6.8600 229.3600 7.7600 ;
      RECT 0.0000 6.5400 230.4600 6.8600 ;
      RECT 1.1000 6.3700 229.3600 6.5400 ;
      RECT 225.2000 5.6400 229.3600 6.3700 ;
      RECT 1.1000 5.6400 5.2600 6.3700 ;
      RECT 225.2000 4.7100 230.4600 5.6400 ;
      RECT 0.0000 4.7100 5.2600 5.6400 ;
      RECT 225.2000 3.8100 229.3600 4.7100 ;
      RECT 1.1000 3.8100 5.2600 4.7100 ;
      RECT 225.2000 3.7700 230.4600 3.8100 ;
      RECT 0.0000 3.7700 5.2600 3.8100 ;
      RECT 0.0000 3.4900 230.4600 3.7700 ;
      RECT 1.1000 3.3700 229.3600 3.4900 ;
      RECT 228.2000 2.5900 229.3600 3.3700 ;
      RECT 1.1000 2.5900 2.2600 3.3700 ;
      RECT 228.2000 0.7700 230.4600 2.5900 ;
      RECT 0.0000 0.7700 2.2600 2.5900 ;
      RECT 0.0000 0.0000 230.4600 0.7700 ;
  END
END S_term_single2

END LIBRARY
