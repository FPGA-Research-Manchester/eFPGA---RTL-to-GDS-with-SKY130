// Copyright 2021 University of Manchester
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//module sky130_v1_wrapper (vddio, vssio, vdda, vssa, vccd, vssd, PAD, clock_pad, Rx_pad, ReceiveLED_pad, s_clk_pad, s_data_pad);
module UoM_eFPGA (vddio, vssio, vdda, vssa, vccd, vssd, PAD, clock_pad, Rx_pad, ReceiveLED_pad, s_clk_pad, s_data_pad, porb_h);

	inout vddio;	// Common 3.3V padframe/ESD power
	inout vssio;	// Common padframe/ESD ground
	inout vdda;	// Management 3.3V power
	inout vssa;	// Common analog ground
	inout vccd;	// Management/Common 1.8V power
	inout vssd;	// Common digital ground

	inout [89:0] PAD;

	input clock_pad;
	// UART configuration port
	input Rx_pad;
	output ReceiveLED_pad;

	// BitBang configuration port
	input s_clk_pad;
	input s_data_pad;

	// Power-up enable
	input porb_h;

	// External USER ports 
	wire [29:0] I_top; 
	wire [29:0] T_top;
	wire [29:0] O_top;

	wire [59:0] OPA;  // go to the CPU
	wire [59:0] OPB;  // go to the CPU
	wire [59:0] RES0; // go to the CPU
	wire [59:0] RES1; // go to the CPU
	wire [59:0] RES2; // go to the CPU
	wire CLK; // This clock can go to the CPU (connects to the fabric LUT wire flops

	// CPU configuration port
	wire SelfWriteStrobe; // must decode address and write enable
	wire [31:0] SelfWriteData; // configuration data write port

	// UART configuration port
	wire Rx;
	wire ComActive;
	wire ReceiveLED;

	// BitBang configuration port
	wire s_clk;
	wire s_data;
	
	wire porb_h;
	
	//simple_por por (
	//	.vdd3v3(vddio),
	//	.vss(vssio),
	//	.porb_h(porb_h)
	//);
	
	eFPGA_top inst_eFPGA_top (
		.I_top(I_top),
		.T_top(T_top),
		.O_top(O_top),
		.OPA(OPA),
		.OPB(OPB),
		.RES0(RES0),
		.RES1(RES1),
		.RES2(RES2),
		.CLK(CLK),
		.SelfWriteStrobe(SelfWriteStrobe),
		.SelfWriteData(SelfWriteData),
		.Rx(Rx),
		.ComActive(ComActive),
		.ReceiveLED(ReceiveLED),
		.s_clk(s_clk),
		.s_data(s_data)
	);

	assign SelfWriteData = RES0[31:0];
	assign SelfWriteStrobe = RES0[32];
	
	//input pads
	wire CLK_loop;
	wire CLK_analog_a,CLK_analog_b;
	wire CLK_vddio_q, CLK_vssio_q;
	sky130_ef_io__gpiov2_pad CLK_in (
		.AMUXBUS_A(CLK_analog_a),
		.AMUXBUS_B(CLK_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(CLK_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(CLK_vssio_q),
		.PAD(clock_pad),
		.OUT(vssd),
		.OE_N(vccd),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(CLK_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		//.INP_DIS(~porb_h), //.INP_DIS(por),
		.INP_DIS(vssd), //for debugging
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vssd, vssd, vccd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(CLK),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(CLK_loop)
	);

	wire Rx_loop;
	wire Rx_analog_a,Rx_analog_b;
	wire Rx_vddio_q, Rx_vssio_q;
	sky130_ef_io__gpiov2_pad Rx_in (
		.AMUXBUS_A(Rx_analog_a),
		.AMUXBUS_B(Rx_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(Rx_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(Rx_vssio_q),
		.PAD(Rx_pad),
		.OUT(vssd),
		.OE_N(vccd),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(Rx_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		//.INP_DIS(~porb_h), //.INP_DIS(por),
		.INP_DIS(vssd), //for debugging
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vssd, vssd, vccd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(Rx),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(Rx_loop)
	);

	wire s_clk_loop;
	wire s_clk_analog_a,s_clk_analog_b;
	wire s_clk_vddio_q, s_clk_vssio_q;
	//sky130_ef_io__gpiov2_pad s_s_clk_in (
	sky130_ef_io__gpiov2_pad s_clk_in (
		.AMUXBUS_A(s_clk_analog_a),
		.AMUXBUS_B(s_clk_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(s_clk_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(s_clk_vssio_q),
		.PAD(s_clk_pad),
		.OUT(vssd),
		.OE_N(vccd),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(s_clk_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		//.INP_DIS(~porb_h), //.INP_DIS(por),
		.INP_DIS(vssd), //for debugging
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vssd, vssd, vccd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(s_clk),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(s_clk_loop)
	);

	wire s_data_loop;
	wire s_data_analog_a,s_data_analog_b;
	wire s_data_vddio_q, s_data_vssio_q;
	sky130_ef_io__gpiov2_pad s_data_in (
		.AMUXBUS_A(s_data_analog_a),
		.AMUXBUS_B(s_data_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(s_data_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(s_data_vssio_q),
		.PAD(s_data_pad),
		.OUT(vssd),
		.OE_N(vccd),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(s_data_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		//.INP_DIS(~porb_h), //.INP_DIS(por),
		.INP_DIS(vssd), //for debugging
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vssd, vssd, vccd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(s_data),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(s_data_loop)
	);

	//output pad
	wire ReceiveLED_loop;
	wire ReceiveLED_analog_a,ReceiveLED_analog_b;
	wire ReceiveLED_vddio_q, ReceiveLED_vssio_q;
	sky130_ef_io__gpiov2_pad ReceiveLED_out (
		.AMUXBUS_A(ReceiveLED_analog_a),
		.AMUXBUS_B(ReceiveLED_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(ReceiveLED_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(ReceiveLED_vssio_q),
		.PAD(ReceiveLED_pad),
		.OUT(ReceiveLED),
		.OE_N(vssd),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(ReceiveLED_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vccd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(ReceiveLED_loop)
	);
	
	//io pads
	wire PAD0_loop;
	wire PAD0_analog_a,PAD0_analog_b;
	wire PAD0_vddio_q, PAD0_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_0 (
		.AMUXBUS_A(PAD0_analog_a),
		.AMUXBUS_B(PAD0_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD0_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD0_vssio_q),
		.PAD(PAD[0]),
		.OUT(I_top[0]),
		.OE_N(T_top[0]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD0_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[0]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD0_loop)
	);

	wire PAD1_loop;
	wire PAD1_analog_a,PAD1_analog_b;
	wire PAD1_vddio_q, PAD1_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_1 (
		.AMUXBUS_A(PAD1_analog_a),
		.AMUXBUS_B(PAD1_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD1_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD1_vssio_q),
		.PAD(PAD[1]),
		.OUT(I_top[1]),
		.OE_N(T_top[1]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD1_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[1]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD1_loop)
	);

	wire PAD2_loop;
	wire PAD2_analog_a,PAD2_analog_b;
	wire PAD2_vddio_q, PAD2_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_2 (
		.AMUXBUS_A(PAD2_analog_a),
		.AMUXBUS_B(PAD2_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD2_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD2_vssio_q),
		.PAD(PAD[2]),
		.OUT(I_top[2]),
		.OE_N(T_top[2]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD2_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[2]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD2_loop)
	);

	wire PAD3_loop;
	wire PAD3_analog_a,PAD3_analog_b;
	wire PAD3_vddio_q, PAD3_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_3 (
		.AMUXBUS_A(PAD3_analog_a),
		.AMUXBUS_B(PAD3_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD3_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD3_vssio_q),
		.PAD(PAD[3]),
		.OUT(I_top[3]),
		.OE_N(T_top[3]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD3_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[3]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD3_loop)
	);

	wire PAD4_loop;
	wire PAD4_analog_a,PAD4_analog_b;
	wire PAD4_vddio_q, PAD4_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_4 (
		.AMUXBUS_A(PAD4_analog_a),
		.AMUXBUS_B(PAD4_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD4_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD4_vssio_q),
		.PAD(PAD[4]),
		.OUT(I_top[4]),
		.OE_N(T_top[4]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD4_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[4]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD4_loop)
	);

	wire PAD5_loop;
	wire PAD5_analog_a,PAD5_analog_b;
	wire PAD5_vddio_q, PAD5_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_5 (
		.AMUXBUS_A(PAD5_analog_a),
		.AMUXBUS_B(PAD5_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD5_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD5_vssio_q),
		.PAD(PAD[5]),
		.OUT(I_top[5]),
		.OE_N(T_top[5]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD5_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[5]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD5_loop)
	);

	wire PAD6_loop;
	wire PAD6_analog_a,PAD6_analog_b;
	wire PAD6_vddio_q, PAD6_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_6 (
		.AMUXBUS_A(PAD6_analog_a),
		.AMUXBUS_B(PAD6_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD6_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD6_vssio_q),
		.PAD(PAD[6]),
		.OUT(I_top[6]),
		.OE_N(T_top[6]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD6_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[6]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD6_loop)
	);

	wire PAD7_loop;
	wire PAD7_analog_a,PAD7_analog_b;
	wire PAD7_vddio_q, PAD7_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_7 (
		.AMUXBUS_A(PAD7_analog_a),
		.AMUXBUS_B(PAD7_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD7_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD7_vssio_q),
		.PAD(PAD[7]),
		.OUT(I_top[7]),
		.OE_N(T_top[7]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD7_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[7]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD7_loop)
	);

	wire PAD8_loop;
	wire PAD8_analog_a,PAD8_analog_b;
	wire PAD8_vddio_q, PAD8_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_8 (
		.AMUXBUS_A(PAD8_analog_a),
		.AMUXBUS_B(PAD8_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD8_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD8_vssio_q),
		.PAD(PAD[8]),
		.OUT(I_top[8]),
		.OE_N(T_top[8]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD8_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[8]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD8_loop)
	);

	wire PAD9_loop;
	wire PAD9_analog_a,PAD9_analog_b;
	wire PAD9_vddio_q, PAD9_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_9 (
		.AMUXBUS_A(PAD9_analog_a),
		.AMUXBUS_B(PAD9_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD9_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD9_vssio_q),
		.PAD(PAD[9]),
		.OUT(I_top[9]),
		.OE_N(T_top[9]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD9_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[9]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD9_loop)
	);

	wire PAD10_loop;
	wire PAD10_analog_a,PAD10_analog_b;
	wire PAD10_vddio_q, PAD10_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_10 (
		.AMUXBUS_A(PAD10_analog_a),
		.AMUXBUS_B(PAD10_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD10_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD10_vssio_q),
		.PAD(PAD[10]),
		.OUT(I_top[10]),
		.OE_N(T_top[10]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD10_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[10]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD10_loop)
	);

	wire PAD11_loop;
	wire PAD11_analog_a,PAD11_analog_b;
	wire PAD11_vddio_q, PAD11_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_11 (
		.AMUXBUS_A(PAD11_analog_a),
		.AMUXBUS_B(PAD11_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD11_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD11_vssio_q),
		.PAD(PAD[11]),
		.OUT(I_top[11]),
		.OE_N(T_top[11]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD11_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[11]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD11_loop)
	);

	wire PAD12_loop;
	wire PAD12_analog_a,PAD12_analog_b;
	wire PAD12_vddio_q, PAD12_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_12 (
		.AMUXBUS_A(PAD12_analog_a),
		.AMUXBUS_B(PAD12_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD12_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD12_vssio_q),
		.PAD(PAD[12]),
		.OUT(I_top[12]),
		.OE_N(T_top[12]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD12_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[12]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD12_loop)
	);

	wire PAD13_loop;
	wire PAD13_analog_a,PAD13_analog_b;
	wire PAD13_vddio_q, PAD13_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_13 (
		.AMUXBUS_A(PAD13_analog_a),
		.AMUXBUS_B(PAD13_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD13_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD13_vssio_q),
		.PAD(PAD[13]),
		.OUT(I_top[13]),
		.OE_N(T_top[13]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD13_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[13]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD13_loop)
	);

	wire PAD14_loop;
	wire PAD14_analog_a,PAD14_analog_b;
	wire PAD14_vddio_q, PAD14_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_14 (
		.AMUXBUS_A(PAD14_analog_a),
		.AMUXBUS_B(PAD14_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD14_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD14_vssio_q),
		.PAD(PAD[14]),
		.OUT(I_top[14]),
		.OE_N(T_top[14]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD14_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[14]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD14_loop)
	);

	wire PAD15_loop;
	wire PAD15_analog_a,PAD15_analog_b;
	wire PAD15_vddio_q, PAD15_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_15 (
		.AMUXBUS_A(PAD15_analog_a),
		.AMUXBUS_B(PAD15_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD15_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD15_vssio_q),
		.PAD(PAD[15]),
		.OUT(I_top[15]),
		.OE_N(T_top[15]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD15_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[15]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD15_loop)
	);

	wire PAD16_loop;
	wire PAD16_analog_a,PAD16_analog_b;
	wire PAD16_vddio_q, PAD16_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_16 (
		.AMUXBUS_A(PAD16_analog_a),
		.AMUXBUS_B(PAD16_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD16_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD16_vssio_q),
		.PAD(PAD[16]),
		.OUT(I_top[16]),
		.OE_N(T_top[16]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD16_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[16]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD16_loop)
	);

	wire PAD17_loop;
	wire PAD17_analog_a,PAD17_analog_b;
	wire PAD17_vddio_q, PAD17_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_17 (
		.AMUXBUS_A(PAD17_analog_a),
		.AMUXBUS_B(PAD17_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD17_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD17_vssio_q),
		.PAD(PAD[17]),
		.OUT(I_top[17]),
		.OE_N(T_top[17]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD17_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[17]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD17_loop)
	);

	wire PAD18_loop;
	wire PAD18_analog_a,PAD18_analog_b;
	wire PAD18_vddio_q, PAD18_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_18 (
		.AMUXBUS_A(PAD18_analog_a),
		.AMUXBUS_B(PAD18_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD18_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD18_vssio_q),
		.PAD(PAD[18]),
		.OUT(I_top[18]),
		.OE_N(T_top[18]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD18_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[18]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD18_loop)
	);

	wire PAD19_loop;
	wire PAD19_analog_a,PAD19_analog_b;
	wire PAD19_vddio_q, PAD19_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_19 (
		.AMUXBUS_A(PAD19_analog_a),
		.AMUXBUS_B(PAD19_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD19_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD19_vssio_q),
		.PAD(PAD[19]),
		.OUT(I_top[19]),
		.OE_N(T_top[19]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD19_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[19]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD19_loop)
	);

	wire PAD20_loop;
	wire PAD20_analog_a,PAD20_analog_b;
	wire PAD20_vddio_q, PAD20_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_20 (
		.AMUXBUS_A(PAD20_analog_a),
		.AMUXBUS_B(PAD20_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD20_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD20_vssio_q),
		.PAD(PAD[20]),
		.OUT(I_top[20]),
		.OE_N(T_top[20]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD20_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[20]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD20_loop)
	);

	wire PAD21_loop;
	wire PAD21_analog_a,PAD21_analog_b;
	wire PAD21_vddio_q, PAD21_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_21 (
		.AMUXBUS_A(PAD21_analog_a),
		.AMUXBUS_B(PAD21_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD21_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD21_vssio_q),
		.PAD(PAD[21]),
		.OUT(I_top[21]),
		.OE_N(T_top[21]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD21_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[21]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD21_loop)
	);

	wire PAD22_loop;
	wire PAD22_analog_a,PAD22_analog_b;
	wire PAD22_vddio_q, PAD22_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_22 (
		.AMUXBUS_A(PAD22_analog_a),
		.AMUXBUS_B(PAD22_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD22_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD22_vssio_q),
		.PAD(PAD[22]),
		.OUT(I_top[22]),
		.OE_N(T_top[22]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD22_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[22]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD22_loop)
	);

	wire PAD23_loop;
	wire PAD23_analog_a,PAD23_analog_b;
	wire PAD23_vddio_q, PAD23_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_23 (
		.AMUXBUS_A(PAD23_analog_a),
		.AMUXBUS_B(PAD23_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD23_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD23_vssio_q),
		.PAD(PAD[23]),
		.OUT(I_top[23]),
		.OE_N(T_top[23]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD23_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[23]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD23_loop)
	);

	wire PAD24_loop;
	wire PAD24_analog_a,PAD24_analog_b;
	wire PAD24_vddio_q, PAD24_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_24 (
		.AMUXBUS_A(PAD24_analog_a),
		.AMUXBUS_B(PAD24_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD24_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD24_vssio_q),
		.PAD(PAD[24]),
		.OUT(I_top[24]),
		.OE_N(T_top[24]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD24_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[24]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD24_loop)
	);

	wire PAD25_loop;
	wire PAD25_analog_a,PAD25_analog_b;
	wire PAD25_vddio_q, PAD25_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_25 (
		.AMUXBUS_A(PAD25_analog_a),
		.AMUXBUS_B(PAD25_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD25_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD25_vssio_q),
		.PAD(PAD[25]),
		.OUT(I_top[25]),
		.OE_N(T_top[25]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD25_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[25]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD25_loop)
	);

	wire PAD26_loop;
	wire PAD26_analog_a,PAD26_analog_b;
	wire PAD26_vddio_q, PAD26_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_26 (
		.AMUXBUS_A(PAD26_analog_a),
		.AMUXBUS_B(PAD26_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD26_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD26_vssio_q),
		.PAD(PAD[26]),
		.OUT(I_top[26]),
		.OE_N(T_top[26]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD26_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[26]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD26_loop)
	);

	wire PAD27_loop;
	wire PAD27_analog_a,PAD27_analog_b;
	wire PAD27_vddio_q, PAD27_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_27 (
		.AMUXBUS_A(PAD27_analog_a),
		.AMUXBUS_B(PAD27_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD27_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD27_vssio_q),
		.PAD(PAD[27]),
		.OUT(I_top[27]),
		.OE_N(T_top[27]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD27_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[27]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD27_loop)
	);

	wire PAD28_loop;
	wire PAD28_analog_a,PAD28_analog_b;
	wire PAD28_vddio_q, PAD28_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_28 (
		.AMUXBUS_A(PAD28_analog_a),
		.AMUXBUS_B(PAD28_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD28_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD28_vssio_q),
		.PAD(PAD[28]),
		.OUT(I_top[28]),
		.OE_N(T_top[28]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD28_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[28]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD28_loop)
	);

	wire PAD29_loop;
	wire PAD29_analog_a,PAD29_analog_b;
	wire PAD29_vddio_q, PAD29_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_29 (
		.AMUXBUS_A(PAD29_analog_a),
		.AMUXBUS_B(PAD29_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD29_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD29_vssio_q),
		.PAD(PAD[29]),
		.OUT(I_top[29]),
		.OE_N(T_top[29]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD29_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(O_top[29]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD29_loop)
	);

	wire PAD30_loop;
	wire PAD30_analog_a,PAD30_analog_b;
	wire PAD30_vddio_q, PAD30_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_30 (
		.AMUXBUS_A(PAD30_analog_a),
		.AMUXBUS_B(PAD30_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD30_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD30_vssio_q),
		.PAD(PAD[30]),
		.OUT(RES1[0]),
		.OE_N(RES2[0]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD30_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[0]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD30_loop)
	);

	wire PAD31_loop;
	wire PAD31_analog_a,PAD31_analog_b;
	wire PAD31_vddio_q, PAD31_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_31 (
		.AMUXBUS_A(PAD31_analog_a),
		.AMUXBUS_B(PAD31_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD31_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD31_vssio_q),
		.PAD(PAD[31]),
		.OUT(RES1[1]),
		.OE_N(RES2[1]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD31_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[1]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD31_loop)
	);

	wire PAD32_loop;
	wire PAD32_analog_a,PAD32_analog_b;
	wire PAD32_vddio_q, PAD32_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_32 (
		.AMUXBUS_A(PAD32_analog_a),
		.AMUXBUS_B(PAD32_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD32_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD32_vssio_q),
		.PAD(PAD[32]),
		.OUT(RES1[2]),
		.OE_N(RES2[2]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD32_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[2]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD32_loop)
	);

	wire PAD33_loop;
	wire PAD33_analog_a,PAD33_analog_b;
	wire PAD33_vddio_q, PAD33_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_33 (
		.AMUXBUS_A(PAD33_analog_a),
		.AMUXBUS_B(PAD33_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD33_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD33_vssio_q),
		.PAD(PAD[33]),
		.OUT(RES1[3]),
		.OE_N(RES2[3]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD33_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[3]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD33_loop)
	);

	wire PAD34_loop;
	wire PAD34_analog_a,PAD34_analog_b;
	wire PAD34_vddio_q, PAD34_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_34 (
		.AMUXBUS_A(PAD34_analog_a),
		.AMUXBUS_B(PAD34_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD34_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD34_vssio_q),
		.PAD(PAD[34]),
		.OUT(RES1[4]),
		.OE_N(RES2[4]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD34_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[4]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD34_loop)
	);

	wire PAD35_loop;
	wire PAD35_analog_a,PAD35_analog_b;
	wire PAD35_vddio_q, PAD35_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_35 (
		.AMUXBUS_A(PAD35_analog_a),
		.AMUXBUS_B(PAD35_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD35_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD35_vssio_q),
		.PAD(PAD[35]),
		.OUT(RES1[5]),
		.OE_N(RES2[5]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD35_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[5]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD35_loop)
	);

	wire PAD36_loop;
	wire PAD36_analog_a,PAD36_analog_b;
	wire PAD36_vddio_q, PAD36_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_36 (
		.AMUXBUS_A(PAD36_analog_a),
		.AMUXBUS_B(PAD36_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD36_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD36_vssio_q),
		.PAD(PAD[36]),
		.OUT(RES1[6]),
		.OE_N(RES2[6]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD36_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[6]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD36_loop)
	);

	wire PAD37_loop;
	wire PAD37_analog_a,PAD37_analog_b;
	wire PAD37_vddio_q, PAD37_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_37 (
		.AMUXBUS_A(PAD37_analog_a),
		.AMUXBUS_B(PAD37_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD37_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD37_vssio_q),
		.PAD(PAD[37]),
		.OUT(RES1[7]),
		.OE_N(RES2[7]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD37_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[7]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD37_loop)
	);

	wire PAD38_loop;
	wire PAD38_analog_a,PAD38_analog_b;
	wire PAD38_vddio_q, PAD38_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_38 (
		.AMUXBUS_A(PAD38_analog_a),
		.AMUXBUS_B(PAD38_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD38_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD38_vssio_q),
		.PAD(PAD[38]),
		.OUT(RES1[8]),
		.OE_N(RES2[8]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD38_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[8]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD38_loop)
	);

	wire PAD39_loop;
	wire PAD39_analog_a,PAD39_analog_b;
	wire PAD39_vddio_q, PAD39_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_39 (
		.AMUXBUS_A(PAD39_analog_a),
		.AMUXBUS_B(PAD39_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD39_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD39_vssio_q),
		.PAD(PAD[39]),
		.OUT(RES1[9]),
		.OE_N(RES2[9]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD39_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[9]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD39_loop)
	);

	wire PAD40_loop;
	wire PAD40_analog_a,PAD40_analog_b;
	wire PAD40_vddio_q, PAD40_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_40 (
		.AMUXBUS_A(PAD40_analog_a),
		.AMUXBUS_B(PAD40_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD40_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD40_vssio_q),
		.PAD(PAD[40]),
		.OUT(RES1[10]),
		.OE_N(RES2[10]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD40_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[10]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD40_loop)
	);

	wire PAD41_loop;
	wire PAD41_analog_a,PAD41_analog_b;
	wire PAD41_vddio_q, PAD41_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_41 (
		.AMUXBUS_A(PAD41_analog_a),
		.AMUXBUS_B(PAD41_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD41_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD41_vssio_q),
		.PAD(PAD[41]),
		.OUT(RES1[11]),
		.OE_N(RES2[11]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD41_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[11]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD41_loop)
	);

	wire PAD42_loop;
	wire PAD42_analog_a,PAD42_analog_b;
	wire PAD42_vddio_q, PAD42_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_42 (
		.AMUXBUS_A(PAD42_analog_a),
		.AMUXBUS_B(PAD42_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD42_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD42_vssio_q),
		.PAD(PAD[42]),
		.OUT(RES1[12]),
		.OE_N(RES2[12]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD42_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[12]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD42_loop)
	);

	wire PAD43_loop;
	wire PAD43_analog_a,PAD43_analog_b;
	wire PAD43_vddio_q, PAD43_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_43 (
		.AMUXBUS_A(PAD43_analog_a),
		.AMUXBUS_B(PAD43_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD43_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD43_vssio_q),
		.PAD(PAD[43]),
		.OUT(RES1[13]),
		.OE_N(RES2[13]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD43_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[13]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD43_loop)
	);

	wire PAD44_loop;
	wire PAD44_analog_a,PAD44_analog_b;
	wire PAD44_vddio_q, PAD44_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_44 (
		.AMUXBUS_A(PAD44_analog_a),
		.AMUXBUS_B(PAD44_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD44_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD44_vssio_q),
		.PAD(PAD[44]),
		.OUT(RES1[14]),
		.OE_N(RES2[14]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD44_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[14]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD44_loop)
	);

	wire PAD45_loop;
	wire PAD45_analog_a,PAD45_analog_b;
	wire PAD45_vddio_q, PAD45_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_45 (
		.AMUXBUS_A(PAD45_analog_a),
		.AMUXBUS_B(PAD45_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD45_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD45_vssio_q),
		.PAD(PAD[45]),
		.OUT(RES1[15]),
		.OE_N(RES2[15]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD45_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[15]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD45_loop)
	);

	wire PAD46_loop;
	wire PAD46_analog_a,PAD46_analog_b;
	wire PAD46_vddio_q, PAD46_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_46 (
		.AMUXBUS_A(PAD46_analog_a),
		.AMUXBUS_B(PAD46_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD46_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD46_vssio_q),
		.PAD(PAD[46]),
		.OUT(RES1[16]),
		.OE_N(RES2[16]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD46_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[16]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD46_loop)
	);

	wire PAD47_loop;
	wire PAD47_analog_a,PAD47_analog_b;
	wire PAD47_vddio_q, PAD47_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_47 (
		.AMUXBUS_A(PAD47_analog_a),
		.AMUXBUS_B(PAD47_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD47_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD47_vssio_q),
		.PAD(PAD[47]),
		.OUT(RES1[17]),
		.OE_N(RES2[17]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD47_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[17]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD47_loop)
	);

	wire PAD48_loop;
	wire PAD48_analog_a,PAD48_analog_b;
	wire PAD48_vddio_q, PAD48_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_48 (
		.AMUXBUS_A(PAD48_analog_a),
		.AMUXBUS_B(PAD48_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD48_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD48_vssio_q),
		.PAD(PAD[48]),
		.OUT(RES1[18]),
		.OE_N(RES2[18]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD48_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[18]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD48_loop)
	);

	wire PAD49_loop;
	wire PAD49_analog_a,PAD49_analog_b;
	wire PAD49_vddio_q, PAD49_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_49 (
		.AMUXBUS_A(PAD49_analog_a),
		.AMUXBUS_B(PAD49_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD49_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD49_vssio_q),
		.PAD(PAD[49]),
		.OUT(RES1[19]),
		.OE_N(RES2[19]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD49_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[19]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD49_loop)
	);

	wire PAD50_loop;
	wire PAD50_analog_a,PAD50_analog_b;
	wire PAD50_vddio_q, PAD50_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_50 (
		.AMUXBUS_A(PAD50_analog_a),
		.AMUXBUS_B(PAD50_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD50_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD50_vssio_q),
		.PAD(PAD[50]),
		.OUT(RES1[20]),
		.OE_N(RES2[20]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD50_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[20]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD50_loop)
	);

	wire PAD51_loop;
	wire PAD51_analog_a,PAD51_analog_b;
	wire PAD51_vddio_q, PAD51_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_51 (
		.AMUXBUS_A(PAD51_analog_a),
		.AMUXBUS_B(PAD51_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD51_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD51_vssio_q),
		.PAD(PAD[51]),
		.OUT(RES1[21]),
		.OE_N(RES2[21]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD51_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[21]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD51_loop)
	);

	wire PAD52_loop;
	wire PAD52_analog_a,PAD52_analog_b;
	wire PAD52_vddio_q, PAD52_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_52 (
		.AMUXBUS_A(PAD52_analog_a),
		.AMUXBUS_B(PAD52_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD52_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD52_vssio_q),
		.PAD(PAD[52]),
		.OUT(RES1[22]),
		.OE_N(RES2[22]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD52_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[22]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD52_loop)
	);

	wire PAD53_loop;
	wire PAD53_analog_a,PAD53_analog_b;
	wire PAD53_vddio_q, PAD53_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_53 (
		.AMUXBUS_A(PAD53_analog_a),
		.AMUXBUS_B(PAD53_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD53_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD53_vssio_q),
		.PAD(PAD[53]),
		.OUT(RES1[23]),
		.OE_N(RES2[23]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD53_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[23]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD53_loop)
	);

	wire PAD54_loop;
	wire PAD54_analog_a,PAD54_analog_b;
	wire PAD54_vddio_q, PAD54_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_54 (
		.AMUXBUS_A(PAD54_analog_a),
		.AMUXBUS_B(PAD54_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD54_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD54_vssio_q),
		.PAD(PAD[54]),
		.OUT(RES1[24]),
		.OE_N(RES2[24]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD54_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[24]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD54_loop)
	);

	wire PAD55_loop;
	wire PAD55_analog_a,PAD55_analog_b;
	wire PAD55_vddio_q, PAD55_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_55 (
		.AMUXBUS_A(PAD55_analog_a),
		.AMUXBUS_B(PAD55_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD55_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD55_vssio_q),
		.PAD(PAD[55]),
		.OUT(RES1[25]),
		.OE_N(RES2[25]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD55_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[25]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD55_loop)
	);

	wire PAD56_loop;
	wire PAD56_analog_a,PAD56_analog_b;
	wire PAD56_vddio_q, PAD56_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_56 (
		.AMUXBUS_A(PAD56_analog_a),
		.AMUXBUS_B(PAD56_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD56_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD56_vssio_q),
		.PAD(PAD[56]),
		.OUT(RES1[26]),
		.OE_N(RES2[26]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD56_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[26]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD56_loop)
	);

	wire PAD57_loop;
	wire PAD57_analog_a,PAD57_analog_b;
	wire PAD57_vddio_q, PAD57_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_57 (
		.AMUXBUS_A(PAD57_analog_a),
		.AMUXBUS_B(PAD57_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD57_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD57_vssio_q),
		.PAD(PAD[57]),
		.OUT(RES1[27]),
		.OE_N(RES2[27]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD57_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[27]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD57_loop)
	);

	wire PAD58_loop;
	wire PAD58_analog_a,PAD58_analog_b;
	wire PAD58_vddio_q, PAD58_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_58 (
		.AMUXBUS_A(PAD58_analog_a),
		.AMUXBUS_B(PAD58_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD58_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD58_vssio_q),
		.PAD(PAD[58]),
		.OUT(RES1[28]),
		.OE_N(RES2[28]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD58_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[28]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD58_loop)
	);

	wire PAD59_loop;
	wire PAD59_analog_a,PAD59_analog_b;
	wire PAD59_vddio_q, PAD59_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_59 (
		.AMUXBUS_A(PAD59_analog_a),
		.AMUXBUS_B(PAD59_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD59_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD59_vssio_q),
		.PAD(PAD[59]),
		.OUT(RES1[29]),
		.OE_N(RES2[29]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD59_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[29]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD59_loop)
	);

	wire PAD60_loop;
	wire PAD60_analog_a,PAD60_analog_b;
	wire PAD60_vddio_q, PAD60_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_60 (
		.AMUXBUS_A(PAD60_analog_a),
		.AMUXBUS_B(PAD60_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD60_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD60_vssio_q),
		.PAD(PAD[60]),
		.OUT(RES1[30]),
		.OE_N(RES2[30]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD60_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[30]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD60_loop)
	);

	wire PAD61_loop;
	wire PAD61_analog_a,PAD61_analog_b;
	wire PAD61_vddio_q, PAD61_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_61 (
		.AMUXBUS_A(PAD61_analog_a),
		.AMUXBUS_B(PAD61_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD61_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD61_vssio_q),
		.PAD(PAD[61]),
		.OUT(RES1[31]),
		.OE_N(RES2[31]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD61_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[31]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD61_loop)
	);

	wire PAD62_loop;
	wire PAD62_analog_a,PAD62_analog_b;
	wire PAD62_vddio_q, PAD62_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_62 (
		.AMUXBUS_A(PAD62_analog_a),
		.AMUXBUS_B(PAD62_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD62_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD62_vssio_q),
		.PAD(PAD[62]),
		.OUT(RES1[32]),
		.OE_N(RES2[32]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD62_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[32]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD62_loop)
	);

	wire PAD63_loop;
	wire PAD63_analog_a,PAD63_analog_b;
	wire PAD63_vddio_q, PAD63_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_63 (
		.AMUXBUS_A(PAD63_analog_a),
		.AMUXBUS_B(PAD63_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD63_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD63_vssio_q),
		.PAD(PAD[63]),
		.OUT(RES1[33]),
		.OE_N(RES2[33]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD63_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[33]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD63_loop)
	);

	wire PAD64_loop;
	wire PAD64_analog_a,PAD64_analog_b;
	wire PAD64_vddio_q, PAD64_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_64 (
		.AMUXBUS_A(PAD64_analog_a),
		.AMUXBUS_B(PAD64_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD64_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD64_vssio_q),
		.PAD(PAD[64]),
		.OUT(RES1[34]),
		.OE_N(RES2[34]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD64_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[34]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD64_loop)
	);

	wire PAD65_loop;
	wire PAD65_analog_a,PAD65_analog_b;
	wire PAD65_vddio_q, PAD65_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_65 (
		.AMUXBUS_A(PAD65_analog_a),
		.AMUXBUS_B(PAD65_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD65_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD65_vssio_q),
		.PAD(PAD[65]),
		.OUT(RES1[35]),
		.OE_N(RES2[35]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD65_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[35]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD65_loop)
	);

	wire PAD66_loop;
	wire PAD66_analog_a,PAD66_analog_b;
	wire PAD66_vddio_q, PAD66_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_66 (
		.AMUXBUS_A(PAD66_analog_a),
		.AMUXBUS_B(PAD66_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD66_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD66_vssio_q),
		.PAD(PAD[66]),
		.OUT(RES1[36]),
		.OE_N(RES2[36]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD66_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[36]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD66_loop)
	);

	wire PAD67_loop;
	wire PAD67_analog_a,PAD67_analog_b;
	wire PAD67_vddio_q, PAD67_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_67 (
		.AMUXBUS_A(PAD67_analog_a),
		.AMUXBUS_B(PAD67_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD67_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD67_vssio_q),
		.PAD(PAD[67]),
		.OUT(RES1[37]),
		.OE_N(RES2[37]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD67_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[37]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD67_loop)
	);

	wire PAD68_loop;
	wire PAD68_analog_a,PAD68_analog_b;
	wire PAD68_vddio_q, PAD68_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_68 (
		.AMUXBUS_A(PAD68_analog_a),
		.AMUXBUS_B(PAD68_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD68_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD68_vssio_q),
		.PAD(PAD[68]),
		.OUT(RES1[38]),
		.OE_N(RES2[38]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD68_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[38]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD68_loop)
	);

	wire PAD69_loop;
	wire PAD69_analog_a,PAD69_analog_b;
	wire PAD69_vddio_q, PAD69_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_69 (
		.AMUXBUS_A(PAD69_analog_a),
		.AMUXBUS_B(PAD69_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD69_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD69_vssio_q),
		.PAD(PAD[69]),
		.OUT(RES1[39]),
		.OE_N(RES2[39]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD69_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[39]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD69_loop)
	);

	wire PAD70_loop;
	wire PAD70_analog_a,PAD70_analog_b;
	wire PAD70_vddio_q, PAD70_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_70 (
		.AMUXBUS_A(PAD70_analog_a),
		.AMUXBUS_B(PAD70_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD70_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD70_vssio_q),
		.PAD(PAD[70]),
		.OUT(RES1[40]),
		.OE_N(RES2[40]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD70_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[40]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD70_loop)
	);

	wire PAD71_loop;
	wire PAD71_analog_a,PAD71_analog_b;
	wire PAD71_vddio_q, PAD71_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_71 (
		.AMUXBUS_A(PAD71_analog_a),
		.AMUXBUS_B(PAD71_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD71_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD71_vssio_q),
		.PAD(PAD[71]),
		.OUT(RES1[41]),
		.OE_N(RES2[41]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD71_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[41]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD71_loop)
	);

	wire PAD72_loop;
	wire PAD72_analog_a,PAD72_analog_b;
	wire PAD72_vddio_q, PAD72_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_72 (
		.AMUXBUS_A(PAD72_analog_a),
		.AMUXBUS_B(PAD72_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD72_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD72_vssio_q),
		.PAD(PAD[72]),
		.OUT(RES1[42]),
		.OE_N(RES2[42]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD72_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[42]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD72_loop)
	);

	wire PAD73_loop;
	wire PAD73_analog_a,PAD73_analog_b;
	wire PAD73_vddio_q, PAD73_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_73 (
		.AMUXBUS_A(PAD73_analog_a),
		.AMUXBUS_B(PAD73_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD73_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD73_vssio_q),
		.PAD(PAD[73]),
		.OUT(RES1[43]),
		.OE_N(RES2[43]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD73_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[43]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD73_loop)
	);

	wire PAD74_loop;
	wire PAD74_analog_a,PAD74_analog_b;
	wire PAD74_vddio_q, PAD74_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_74 (
		.AMUXBUS_A(PAD74_analog_a),
		.AMUXBUS_B(PAD74_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD74_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD74_vssio_q),
		.PAD(PAD[74]),
		.OUT(RES1[44]),
		.OE_N(RES2[44]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD74_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[44]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD74_loop)
	);

	wire PAD75_loop;
	wire PAD75_analog_a,PAD75_analog_b;
	wire PAD75_vddio_q, PAD75_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_75 (
		.AMUXBUS_A(PAD75_analog_a),
		.AMUXBUS_B(PAD75_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD75_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD75_vssio_q),
		.PAD(PAD[75]),
		.OUT(RES1[45]),
		.OE_N(RES2[45]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD75_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[45]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD75_loop)
	);

	wire PAD76_loop;
	wire PAD76_analog_a,PAD76_analog_b;
	wire PAD76_vddio_q, PAD76_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_76 (
		.AMUXBUS_A(PAD76_analog_a),
		.AMUXBUS_B(PAD76_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD76_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD76_vssio_q),
		.PAD(PAD[76]),
		.OUT(RES1[46]),
		.OE_N(RES2[46]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD76_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[46]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD76_loop)
	);

	wire PAD77_loop;
	wire PAD77_analog_a,PAD77_analog_b;
	wire PAD77_vddio_q, PAD77_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_77 (
		.AMUXBUS_A(PAD77_analog_a),
		.AMUXBUS_B(PAD77_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD77_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD77_vssio_q),
		.PAD(PAD[77]),
		.OUT(RES1[47]),
		.OE_N(RES2[47]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD77_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[47]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD77_loop)
	);

	wire PAD78_loop;
	wire PAD78_analog_a,PAD78_analog_b;
	wire PAD78_vddio_q, PAD78_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_78 (
		.AMUXBUS_A(PAD78_analog_a),
		.AMUXBUS_B(PAD78_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD78_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD78_vssio_q),
		.PAD(PAD[78]),
		.OUT(RES1[48]),
		.OE_N(RES2[48]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD78_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[48]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD78_loop)
	);

	wire PAD79_loop;
	wire PAD79_analog_a,PAD79_analog_b;
	wire PAD79_vddio_q, PAD79_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_79 (
		.AMUXBUS_A(PAD79_analog_a),
		.AMUXBUS_B(PAD79_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD79_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD79_vssio_q),
		.PAD(PAD[79]),
		.OUT(RES1[49]),
		.OE_N(RES2[49]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD79_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[49]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD79_loop)
	);

	wire PAD80_loop;
	wire PAD80_analog_a,PAD80_analog_b;
	wire PAD80_vddio_q, PAD80_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_80 (
		.AMUXBUS_A(PAD80_analog_a),
		.AMUXBUS_B(PAD80_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD80_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD80_vssio_q),
		.PAD(PAD[80]),
		.OUT(RES1[50]),
		.OE_N(RES2[50]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD80_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[50]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD80_loop)
	);

	wire PAD81_loop;
	wire PAD81_analog_a,PAD81_analog_b;
	wire PAD81_vddio_q, PAD81_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_81 (
		.AMUXBUS_A(PAD81_analog_a),
		.AMUXBUS_B(PAD81_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD81_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD81_vssio_q),
		.PAD(PAD[81]),
		.OUT(RES1[51]),
		.OE_N(RES2[51]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD81_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[51]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD81_loop)
	);

	wire PAD82_loop;
	wire PAD82_analog_a,PAD82_analog_b;
	wire PAD82_vddio_q, PAD82_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_82 (
		.AMUXBUS_A(PAD82_analog_a),
		.AMUXBUS_B(PAD82_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD82_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD82_vssio_q),
		.PAD(PAD[82]),
		.OUT(RES1[52]),
		.OE_N(RES2[52]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD82_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[52]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD82_loop)
	);

	wire PAD83_loop;
	wire PAD83_analog_a,PAD83_analog_b;
	wire PAD83_vddio_q, PAD83_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_83 (
		.AMUXBUS_A(PAD83_analog_a),
		.AMUXBUS_B(PAD83_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD83_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD83_vssio_q),
		.PAD(PAD[83]),
		.OUT(RES1[53]),
		.OE_N(RES2[53]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD83_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[53]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD83_loop)
	);

	wire PAD84_loop;
	wire PAD84_analog_a,PAD84_analog_b;
	wire PAD84_vddio_q, PAD84_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_84 (
		.AMUXBUS_A(PAD84_analog_a),
		.AMUXBUS_B(PAD84_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD84_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD84_vssio_q),
		.PAD(PAD[84]),
		.OUT(RES1[54]),
		.OE_N(RES2[54]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD84_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[54]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD84_loop)
	);

	wire PAD85_loop;
	wire PAD85_analog_a,PAD85_analog_b;
	wire PAD85_vddio_q, PAD85_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_85 (
		.AMUXBUS_A(PAD85_analog_a),
		.AMUXBUS_B(PAD85_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD85_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD85_vssio_q),
		.PAD(PAD[85]),
		.OUT(RES1[55]),
		.OE_N(RES2[55]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD85_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[55]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD85_loop)
	);

	wire PAD86_loop;
	wire PAD86_analog_a,PAD86_analog_b;
	wire PAD86_vddio_q, PAD86_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_86 (
		.AMUXBUS_A(PAD86_analog_a),
		.AMUXBUS_B(PAD86_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD86_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD86_vssio_q),
		.PAD(PAD[86]),
		.OUT(RES1[56]),
		.OE_N(RES2[56]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD86_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[56]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD86_loop)
	);

	wire PAD87_loop;
	wire PAD87_analog_a,PAD87_analog_b;
	wire PAD87_vddio_q, PAD87_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_87 (
		.AMUXBUS_A(PAD87_analog_a),
		.AMUXBUS_B(PAD87_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD87_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD87_vssio_q),
		.PAD(PAD[87]),
		.OUT(RES1[57]),
		.OE_N(RES2[57]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD87_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[57]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD87_loop)
	);

	wire PAD88_loop;
	wire PAD88_analog_a,PAD88_analog_b;
	wire PAD88_vddio_q, PAD88_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_88 (
		.AMUXBUS_A(PAD88_analog_a),
		.AMUXBUS_B(PAD88_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD88_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD88_vssio_q),
		.PAD(PAD[88]),
		.OUT(RES1[58]),
		.OE_N(RES2[58]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD88_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[58]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD88_loop)
	);

	wire PAD89_loop;
	wire PAD89_analog_a,PAD89_analog_b;
	wire PAD89_vddio_q, PAD89_vssio_q;
	sky130_ef_io__gpiov2_pad inst_io_89 (
		.AMUXBUS_A(PAD89_analog_a),
		.AMUXBUS_B(PAD89_analog_b),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(PAD89_vddio_q),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q(PAD89_vssio_q),
		.PAD(PAD[89]),
		.OUT(RES1[59]),
		.OE_N(RES2[59]),
		.HLD_H_N(vddio),
		.ENABLE_H(porb_h),
		.ENABLE_INP_H(PAD89_loop),
		.ENABLE_VDDA_H(porb_h),
		.ENABLE_VSWITCH_H(vssa),
		.ENABLE_VDDIO(vccd),
		.INP_DIS(vssd), //.INP_DIS(INPUT_DIS),
		.IB_MODE_SEL(vssd),
		.VTRIP_SEL(vssd),
		.SLOW(vssd),
		.HLD_OVR(vssd),
		.ANALOG_EN(vssd),
		.ANALOG_SEL(vssd),
		.ANALOG_POL(vssd),
		.DM({vccd, vccd, vssd}),
		.PAD_A_NOESD_H(),
		.PAD_A_ESD_0_H(),
		.PAD_A_ESD_1_H(),
		.IN(OPA[59]),
		.IN_H(),
		.TIE_HI_ESD(),
		.TIE_LO_ESD(PAD89_loop)
	);

	//Power pads
	sky130_ef_io__vccd_lvc_pad pad_vccd_l (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vccd_lvc_pad pad_vccd_t (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vccd_lvc_pad pad_vccd_r (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vccd_lvc_pad pad_vccd_b (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssd_lvc_pad pad_vssd_l (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssd_lvc_pad pad_vssd_t (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssd_lvc_pad pad_vssd_r (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssd_lvc_pad pad_vssd_b (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vddio_lvc_pad pad_vddio_t (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssio_lvc_pad pad_vssio_t (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vddio_lvc_pad pad_vddio_b (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssio_lvc_pad pad_vssio_b (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vdda_lvc_pad pad_vdda_t (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssa_lvc_pad pad_vssa_t (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vdda_lvc_pad pad_vdda_b (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

	sky130_ef_io__vssa_lvc_pad pad_vssa_b (
		.AMUXBUS_A(),
		.AMUXBUS_B(),
		.DRN_LVC1(),
		.DRN_LVC2(),
		.SRC_BDY_LVC1(),
		.SRC_BDY_LVC2(),
		.BDY2_B2B(),
		.VSSA(vssa),
		.VDDA(vdda),
		.VSWITCH(vddio),
		.VDDIO_Q(),
		.VCCHIB(vccd),
		.VDDIO(vddio),
		.VCCD(vccd),
		.VSSIO(vssio),
		.VSSD(vssd),
		.VSSIO_Q()
		);

endmodule



