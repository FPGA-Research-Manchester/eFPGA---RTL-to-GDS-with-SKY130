##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Thu Apr 22 17:29:07 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RegFile
  CLASS BLOCK ;
  SIZE 230.4600 BY 229.8400 ;
  FOREIGN RegFile 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5652 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.752 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 229.5100 19.1750 229.8400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.2995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.653 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.3658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.088 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 229.5100 17.7950 229.8400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.87725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.385 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.7628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.6208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.448 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 229.5100 16.4150 229.8400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.68685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.787 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.8188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.504 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 229.5100 15.4950 229.8400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.56825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.845 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 28.5538 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 142.695 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 29.5850 229.5100 29.7550 229.8400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.888 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 229.5100 28.3750 229.8400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.22445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.1646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 229.5100 26.9950 229.8400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 73.0625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.65 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 229.5100 26.0750 229.8400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.8278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 229.5100 24.6950 229.8400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.5992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.922 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 23.1450 229.5100 23.3150 229.8400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.226 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 229.5100 21.9350 229.8400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.7428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.3850 229.5100 20.5550 229.8400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.2226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 338.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 40.1650 229.5100 40.3350 229.8400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.5394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 340.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 229.5100 38.9550 229.8400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.4958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 344.448 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 37.8650 229.5100 38.0350 229.8400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2424 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.245 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.2148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 337.616 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 229.5100 36.6550 229.8400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.6126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.208 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.1050 229.5100 35.2750 229.8400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.38005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.153 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5212 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.757 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.0298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 299.296 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.7250 229.5100 33.8950 229.8400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.84245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.697 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.2868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 306 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 229.5100 32.5150 229.8400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.0286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 315.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.9650 229.5100 31.1350 229.8400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.0732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.248 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 229.5100 61.9550 229.8400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.18405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1618 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7315 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.1184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.474 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 229.5100 60.5750 229.8400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.1528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.952 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.0250 229.5100 59.1950 229.8400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.3968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 229.5100 57.8150 229.8400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.9425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.3068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.44 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 229.5100 56.4350 229.8400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.53045 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.977 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.36 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 229.5100 55.0550 229.8400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 229.5100 53.6750 229.8400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.05065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.589 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.937 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 229.5100 52.2950 229.8400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.05105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.1986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 229.5100 50.9150 229.8400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.318 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.516 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 49.8250 229.5100 49.9950 229.8400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.369 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 183.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.2116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 48.4450 229.5100 48.6150 229.8400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.438 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 229.5100 47.2350 229.8400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.366 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 229.5100 45.8550 229.8400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.07105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.613 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.7368 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.647 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 44.3050 229.5100 44.4750 229.8400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.68385 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.981 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 22.5324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 112.585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.0668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 229.5100 43.0950 229.8400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.16365 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.369 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 24.5624 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 122.735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.776 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 229.5100 41.7150 229.8400 ;
    END
  END N4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.5555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.8506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 117.039 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 604.216 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.765437 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 0.0000 19.1750 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.8908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8775 LAYER met4  ;
    ANTENNAMAXAREACAR 124.276 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 642.081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.770981 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 0.0000 17.7950 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.95245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.297 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.0105 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 117.511 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 598.451 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.804762 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 0.0000 16.4150 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.99325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.002 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.4016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 76.2382 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 371.018 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.275017 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.95245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.297 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.0668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.16 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7325 LAYER met3  ;
    ANTENNAMAXAREACAR 35.2498 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 180.099 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.230765 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 29.5850 0.0000 29.7550 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.95245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.297 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.757 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 30.0562 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 148.228 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.379394 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 0.0000 28.3750 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.462 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7325 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7726 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.1434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.246522 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 0.0000 26.9950 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.6348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.83 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met2  ;
    ANTENNAMAXAREACAR 9.33441 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.1663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 0.0000 26.0750 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.1912 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 70.8785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7325 LAYER met2  ;
    ANTENNAMAXAREACAR 8.55224 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.4687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.246522 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 0.0000 24.6950 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.33705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.573 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.4016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.1228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met3  ;
    ANTENNAMAXAREACAR 14.7148 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.0024 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.174007 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 23.1450 0.0000 23.3150 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.19625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.551 LAYER li1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER li1  ;
    ANTENNAMAXAREACAR 2.95791 LAYER li1  ;
    ANTENNAMAXSIDEAREACAR 3.43569 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 3.06997 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 3.98249 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    ANTENNAGATEAREA 1.7325 LAYER met2  ;
    ANTENNAMAXAREACAR 9.68993 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.8212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 0.0000 21.9350 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.5523 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.583 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met1  ;
    ANTENNAMAXAREACAR 20.9367 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 61.7542 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.233535 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 20.3850 0.0000 20.5550 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22145 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.437 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.5124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.4845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.3886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 79.1265 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 349.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.974603 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 40.1650 0.0000 40.3350 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.7058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 105.824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 525.773 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.26147 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 0.0000 38.9550 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 59.3316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 90.0873 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 436.597 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.488017 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 37.8650 0.0000 38.0350 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.8108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 227.036 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 0.0000 36.6550 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.7718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 35.1625 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.609 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.316364 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 35.1050 0.0000 35.2750 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.3378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6536 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.017 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.272323 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 33.7250 0.0000 33.8950 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.8888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.116 LAYER met4  ;
    ANTENNAMAXAREACAR 38.8757 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.026 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.337282 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 0.0000 32.5150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.0418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 61.7874 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.137 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.401616 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 30.9650 0.0000 31.1350 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.7288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 49.1036 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 252.839 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 0.0000 61.9550 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.5468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.72 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 53.6369 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 264.909 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 0.0000 60.5750 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 22.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.541 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.7068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.1848 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.299 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 59.0250 0.0000 59.1950 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.846 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.818 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.28121 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.0114 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 0.0000 57.8150 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.7576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.364 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.466 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.98774 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.4667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 85.4509 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 453.451 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 0.0000 55.0550 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.8076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 103.964 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 28.32 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 140.369 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 0.0000 53.6750 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.9072 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.9172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.598 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 23.0943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.301 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7507 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.868 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 0.0000 50.9150 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.8556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 139.16 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 42.3519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 202.845 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 49.8250 0.0000 49.9950 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 51.3712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 48.4450 0.0000 48.6150 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.2508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 225.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 58.9618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 312.944 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 0.0000 47.2350 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.87465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.029 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 22.9747 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.283 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.316364 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 0.0000 45.8550 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.1858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 29.9747 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.342 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.272323 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 44.3050 0.0000 44.4750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3635 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6295 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.779 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.455038 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 0.0000 43.0950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.93505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.453 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.8718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1161 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 186.329 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 0.0000 41.7150 0.3300 ;
    END
  END N4END[0]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 67.4200 230.4600 67.5600 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.3846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 338.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 66.0600 230.4600 66.2000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.851 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.4888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 64.7000 230.4600 64.8400 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.4318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.44 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 63.0000 230.4600 63.1400 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 79.6600 230.4600 79.8000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 77.9600 230.4600 78.1000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 76.6000 230.4600 76.7400 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 75.2400 230.4600 75.3800 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 224.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 73.5400 230.4600 73.6800 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.88 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.4148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 72.1800 230.4600 72.3200 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.72 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.2566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 70.4800 230.4600 70.6200 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.605 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 302.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.6218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 69.1200 230.4600 69.2600 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.686 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 91.5600 230.4600 91.7000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.0902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.225 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 90.2000 230.4600 90.3400 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.651 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.3798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.496 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 88.5000 230.4600 88.6400 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 87.1400 230.4600 87.2800 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.5988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.664 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 85.7800 230.4600 85.9200 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 84.0800 230.4600 84.2200 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.5694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 82.7200 230.4600 82.8600 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.993 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.6628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 81.0200 230.4600 81.1600 ;
    END
  END E2BEGb[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.7428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.432 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 109.5800 230.4600 109.7200 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 108.2200 230.4600 108.3600 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 106.8600 230.4600 107.0000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 105.1600 230.4600 105.3000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.2318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.933 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 103.8000 230.4600 103.9400 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 102.1000 230.4600 102.2400 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 100.7400 230.4600 100.8800 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.2048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 99.0400 230.4600 99.1800 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 97.6800 230.4600 97.8200 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 96.3200 230.4600 96.4600 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.211 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.8218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 94.6200 230.4600 94.7600 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 93.2600 230.4600 93.4000 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2975 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1295 LAYER met4  ;
    ANTENNAMAXAREACAR 105.149 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 507.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.4200 0.4850 67.5600 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.96 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.99 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.0126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.377 LAYER met4  ;
    ANTENNAMAXAREACAR 61.9031 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.02 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.692328 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.0600 0.4850 66.2000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.8498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 83.2855 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.587 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.606707 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.7000 0.4850 64.8400 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.3794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 74.1653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.598 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.396229 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 63.0000 0.4850 63.1400 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.98 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 304.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.7458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 15.9139 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.4133 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 79.6600 0.4850 79.8000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 263.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 10.743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 43.0391 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.302559 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.9600 0.4850 78.1000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.5488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 18.374 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.7135 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.167273 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 76.6000 0.4850 76.7400 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.1404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 15.2994 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 72.7559 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.231246 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.2400 0.4850 75.3800 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.653 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 222.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.3428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 14.0981 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 71.5572 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.106182 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.5400 0.4850 73.6800 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 44.0293 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 222.949 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.352458 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 72.1800 0.4850 72.3200 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 8.78483 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.5919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0960269 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.4800 0.4850 70.6200 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.481 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.6576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 13.1964 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.2896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.185791 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 69.1200 0.4850 69.2600 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.6246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 58.9102 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.479 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.368969 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.5600 0.4850 91.7000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.1468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5277 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.209 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.895953 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.2000 0.4850 90.3400 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.6396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 51.5975 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.43 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.555072 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.5000 0.4850 88.6400 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.2885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.7028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 38.9259 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.744 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.461484 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.1400 0.4850 87.2800 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.2275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5325 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.5165 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.7800 0.4850 85.9200 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.3448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.976 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 50.4427 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 254.76 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.261549 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.0800 0.4850 84.2200 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1049 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.1766 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.7200 0.4850 82.8600 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 16.4119 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.096 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.0200 0.4850 81.1600 ;
    END
  END E2END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 293.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.5188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.7316 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.824 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.5800 0.4850 109.7200 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.76539 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.2929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.2200 0.4850 108.3600 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 39.2296 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 190.253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.7631 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.3845 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.1600 0.4850 105.3000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.904 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.979 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.2126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.1833 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.858 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1428 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.7394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.1000 0.4850 102.2400 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.309 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.2028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.5879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.252 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.7400 0.4850 100.8800 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 44.3389 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.899 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.0400 0.4850 99.1800 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.23704 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.9946 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.6800 0.4850 97.8200 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2653 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.523 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.5844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 30.8652 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.926 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.3200 0.4850 96.4600 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.844 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 32.9396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.6200 0.4850 94.7600 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.5878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 30.0088 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 138.726 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.455758 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.2600 0.4850 93.4000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.47005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.553 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.4 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.646 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 0.0000 65.6350 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.6732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.816 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 0.0000 64.2550 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.76165 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.249 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.35705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.773 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.1788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.424 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.0050 0.0000 88.1750 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.64605 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.113 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.6778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 86.6250 0.0000 86.7950 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.64605 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.113 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.8504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 0.0000 85.8750 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.9708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 325.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 0.0000 84.4950 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.8408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.086 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 0.0000 83.1150 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.9798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 293.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 0.0000 81.7350 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.7236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 324.8 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 0.0000 80.3550 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0972 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.284 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 78.8050 0.0000 78.9750 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.0008 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.9265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 0.0000 77.5950 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.4385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 76.0450 0.0000 76.2150 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER li1  ;
    ANTENNAPARTIALMETALAREA 4.31035 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5 LAYER li1  ;
    PORT
      LAYER li1 ;
        RECT 74.6650 0.0000 74.8350 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.4652 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.289 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 0.0000 73.9150 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.1168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.51 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.5508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.68 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.11 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.4725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.178 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 0.0000 69.7750 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9028 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.477 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 0.0000 68.3950 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.347 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 109.6250 0.0000 109.7950 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1601 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.2866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.136 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.2450 0.0000 108.4150 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.825 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.2976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.528 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 106.8650 0.0000 107.0350 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.2234 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.6778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.4850 0.0000 105.6550 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.2076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 75.9605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.034 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 104.1050 0.0000 104.2750 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.7846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 319.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.7250 0.0000 102.8950 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.1976 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.9105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.65 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 101.3450 0.0000 101.5150 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 16.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.088 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9650 0.0000 100.1350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.805 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 15.965 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.751 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 98.5850 0.0000 98.7550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 15.9996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.961 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 97.6650 0.0000 97.8350 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.1344 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 306.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 96.2850 0.0000 96.4550 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.5866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 94.9050 0.0000 95.0750 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 17.1252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.589 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 93.5250 0.0000 93.6950 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.31965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.729 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2296 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.6028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.352 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.1450 0.0000 92.3150 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.5126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.008 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 90.7650 0.0000 90.9350 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.3108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 89.3850 0.0000 89.5550 0.3300 ;
    END
  END S4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3144 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.768 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met2  ;
    ANTENNAMAXAREACAR 34.8238 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.693 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.518971 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 229.5100 67.0150 229.8400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.6148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 39.4813 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 196.132 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.777444 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 229.5100 65.6350 229.8400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.8016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met3  ;
    ANTENNAMAXAREACAR 39.5372 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 176.94 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.626066 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 229.5100 64.2550 229.8400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.7128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 97.2446 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 508.406 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530928 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 229.5100 62.8750 229.8400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.4056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 46.1555 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.163 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.141212 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 88.0050 229.5100 88.1750 229.8400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3268 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.5565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.2938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 39.3074 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 206.735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 86.6250 229.5100 86.7950 229.8400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.58825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.045 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.6488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 44.3278 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.426 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.141212 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 229.5100 85.8750 229.8400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.3096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 53.4569 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 229.5100 84.4950 229.8400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0536 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1535 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.6768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 46.887 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.78 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.141212 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 229.5100 83.1150 229.8400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.35705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.773 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.3146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 34.1737 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.684 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.200943 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 229.5100 81.7350 229.8400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 61.9566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 52.9772 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 279.213 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.106182 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 229.5100 80.3550 229.8400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 64.8456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 346.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3521 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.821 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.141212 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 78.8050 229.5100 78.9750 229.8400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.0926 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.3855 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.1524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.644 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2228 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.1202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 229.5100 77.5950 229.8400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.58825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.045 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.0756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 82.8986 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 439.089 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 76.0450 229.5100 76.2150 229.8400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.246 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0887 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.2204 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.259486 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 74.6650 229.5100 74.8350 229.8400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.79 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.0535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 229.5100 73.9150 229.8400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.954 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1123 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.8505 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 229.5100 72.5350 229.8400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.15354 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.5 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 229.5100 71.1550 229.8400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.6168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4916 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.099 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423165 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 229.5100 69.7750 229.8400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.3598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 95.3138 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 461.254 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.746967 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 229.5100 68.3950 229.8400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.6452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 68.1485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.6748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.7046 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.373 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 109.6250 229.5100 109.7950 229.8400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.232 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.0825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.70707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.5455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 108.2450 229.5100 108.4150 229.8400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5364 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.6045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.6598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.9228 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.867 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 106.8650 229.5100 107.0350 229.8400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.0928 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 75.3865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.2848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.1174 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.525 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 105.4850 229.5100 105.6550 229.8400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.2244 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.0445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 290.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.8831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.51 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 104.1050 229.5100 104.2750 229.8400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.1465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.327 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.4768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8813 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.459 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 102.7250 229.5100 102.8950 229.8400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.75905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.893 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.2932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.392 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 15.506 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 76.299 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 101.3450 229.5100 101.5150 229.8400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.198 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.9125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.53051 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.2242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 99.9650 229.5100 100.1350 229.8400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.612 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.7598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 93.4035 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 493.896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 98.5850 229.5100 98.7550 229.8400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.41225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.8828 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.3365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.368 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.63434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.7771 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 97.6650 229.5100 97.8350 229.8400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22145 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.437 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.9064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 59.458 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 16.3319 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 80.4283 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 96.2850 229.5100 96.4550 229.8400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.643 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 14.273 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 59.67 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 94.9050 229.5100 95.0750 229.8400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1432 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.679 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 19.5325 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 78.1192 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0583838 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 93.5250 229.5100 93.6950 229.8400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.47015 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.891 LAYER li1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER li1  ;
    ANTENNAMAXAREACAR 4.9902 LAYER li1  ;
    ANTENNAMAXSIDEAREACAR 5.8404 LAYER li1  ;
    PORT
      LAYER li1 ;
        RECT 92.1450 229.5100 92.3150 229.8400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.3325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 65.3311 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 347.527 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 90.7650 229.5100 90.9350 229.8400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.9816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.79 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2428 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.696 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 89.3850 229.5100 89.5550 229.8400 ;
    END
  END S4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.176 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.4800 0.4850 19.6200 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.7800 0.4850 17.9200 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.4200 0.4850 16.5600 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.0600 0.4850 15.2000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.1008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.3800 0.4850 31.5200 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.5168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.0200 0.4850 30.1600 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.3200 0.4850 28.4600 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.5424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 26.9600 0.4850 27.1000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.544 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.6000 0.4850 25.7400 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.9758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.9000 0.4850 24.0400 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.0298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 315.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.9728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.1138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.744 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 45.4218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.9200 0.4850 42.0600 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.4678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.632 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.708 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.0518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 198.08 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.8600 0.4850 39.0000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.5000 0.4850 37.6400 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.4478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.1400 0.4850 36.2800 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.4400 0.4850 34.5800 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.8578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.0800 0.4850 33.2200 ;
    END
  END W2BEGb[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.8938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.6400 0.4850 61.7800 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.092 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.029 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.5800 0.4850 58.7200 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 57.2200 0.4850 57.3600 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.6884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.5200 0.4850 55.6600 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 60.6498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 323.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 54.1600 0.4850 54.3000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.4600 0.4850 52.6000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.017 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.3618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 338.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.1000 0.4850 51.2400 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.0778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.4000 0.4850 49.5400 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.4838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.0400 0.4850 48.1800 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.223 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.9800 0.4850 45.1200 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.261 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.3676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 55.2957 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.167 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 19.4800 230.4600 19.6200 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.324 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.4306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 52.8824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 270.595 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.366581 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 17.7800 230.4600 17.9200 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.2108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 65.9482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.541258 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 16.4200 230.4600 16.5600 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 31.6516 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 146.706 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.4265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.344 LAYER met3  ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 70.3465 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 340.913 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.08308 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 71.3262 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.08308 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 15.0600 230.4600 15.2000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.491 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 3.71036 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.4419 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0765657 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 31.3800 230.4600 31.5200 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.4478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 15.8335 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.7786 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0738586 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 30.0200 230.4600 30.1600 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.1378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 235.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 39.0802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 199.656 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.108889 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 28.3200 230.4600 28.4600 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.6548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 25.9633 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 125.686 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.167273 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 26.9600 230.4600 27.1000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 26.2642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.106182 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 25.6000 230.4600 25.7400 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.7618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7716 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.464 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.136162 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 23.9000 230.4600 24.0400 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 60.5148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 323.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 50.9223 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 268.924 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.136162 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 22.5400 230.4600 22.6800 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.4468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0673 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.945 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0738586 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 20.8400 230.4600 20.9800 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.03556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.0697 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 43.6200 230.4600 43.7600 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0339 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.8535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 41.9200 230.4600 42.0600 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.4416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 62.8412 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 329.444 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 40.5600 230.4600 40.7000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.9076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 81.1412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 432.489 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 38.8600 230.4600 39.0000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 106.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.7058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 255.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 11.6481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.4808 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 37.5000 230.4600 37.6400 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.2564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 12.8281 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 66.8747 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 36.1400 230.4600 36.2800 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.5416 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 66.797 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.868 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 34.4400 230.4600 34.5800 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.9048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 35.0188 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 182.806 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 33.0800 230.4600 33.2200 ;
    END
  END W2END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.8766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.4574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 360.078 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 61.6400 230.4600 61.7800 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.2932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.5906 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.353 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 59.9400 230.4600 60.0800 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.30168 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.0774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 58.5800 230.4600 58.7200 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.9103 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.6586 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 57.2200 230.4600 57.3600 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.9856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.0539 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 336.11 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 55.5200 230.4600 55.6600 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.12754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.1886 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 54.1600 230.4600 54.3000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.8786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.6269 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 371.18 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 52.4600 230.4600 52.6000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.6384 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.6353 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.113 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 51.1000 230.4600 51.2400 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.79825 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.503 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 49.4000 230.4600 49.5400 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.8286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 96.1876 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 511.763 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 48.0400 230.4600 48.1800 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.1768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.2424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 44.2861 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 237.691 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 46.6800 230.4600 46.8200 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.4596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 41.4594 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 44.9800 230.4600 45.1200 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9264 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 7.26502 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 37.8865 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 114.3900 0.0000 114.6900 0.8000 ;
    END
  END UserCLK
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met2  ;
    ANTENNAMAXAREACAR 18.325 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.5963 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.63957 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 48.3799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 225.913 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.63957 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 214.3000 0.4850 214.4400 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.7466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6965 LAYER met4  ;
    ANTENNAMAXAREACAR 90.4412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 466.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 211.5800 0.4850 211.7200 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.699 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.0292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 55.099 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.832 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.983016 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 208.5200 0.4850 208.6600 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 40.3674 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.609 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674318 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 205.4600 0.4850 205.6000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.9103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 22.7409 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 84.3113 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.493006 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.8516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.816 LAYER met4  ;
    ANTENNAGATEAREA 1.5375 LAYER met4  ;
    ANTENNAMAXAREACAR 43.3252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.607 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.4000 0.4850 202.5400 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.5923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 37.1159 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 186.797 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.481076 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.9207 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.376 LAYER met4  ;
    ANTENNAGATEAREA 1.6965 LAYER met4  ;
    ANTENNAMAXAREACAR 72.4174 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.393 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 199.3400 0.4850 199.4800 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.0928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met3  ;
    ANTENNAMAXAREACAR 45.6584 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 204.419 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.798679 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 196.2800 0.4850 196.4200 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.5903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 52.5917 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.659 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.622956 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.1765 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.544 LAYER met4  ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 62.7355 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.008 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.2200 0.4850 193.3600 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 9.34079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.2929 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.360988 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.1193 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.568 LAYER met3  ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 27.3046 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.924 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.21529 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.2916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.496 LAYER met4  ;
    ANTENNAGATEAREA 1.5375 LAYER met4  ;
    ANTENNAMAXAREACAR 80.6306 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.211 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.21529 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.1600 0.4850 190.3000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 5.84124 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8516 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.261912 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.1018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.48 LAYER met3  ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 58.6229 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 260.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.6798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.096 LAYER met4  ;
    ANTENNAGATEAREA 1.6965 LAYER met4  ;
    ANTENNAMAXAREACAR 76.7071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.214 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2504 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 187.1000 0.4850 187.2400 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.598 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6981 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.8711 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.0983 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.064 LAYER met3  ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 71.2998 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 358.914 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.2 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.24 LAYER met4  ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 73.8789 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.795 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 184.0400 0.4850 184.1800 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 26.8758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.653 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.827358 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.0276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.888 LAYER met3  ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1306 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.449 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.877673 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3015 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.544 LAYER met4  ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 66.1964 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 331.382 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.877673 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 180.9800 0.4850 181.1200 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 193.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.0497 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met4  ;
    ANTENNAMAXAREACAR 34.8412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 142.995 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.37673 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.9200 0.4850 178.0600 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.0977 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6965 LAYER met4  ;
    ANTENNAMAXAREACAR 35.4762 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.686 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.407128 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.8600 0.4850 175.0000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.21 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.9135 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 42.9771 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.969 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.651782 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 171.8000 0.4850 171.9400 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.5738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 46.2514 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.81 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.667798 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 168.7400 0.4850 168.8800 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.957 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.9288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 46.5927 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 233.252 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.6800 0.4850 165.8200 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 42.224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.731 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381305 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 162.6200 0.4850 162.7600 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.2563 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 69.9888 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.713 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666038 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 159.5600 0.4850 159.7000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 58.996 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 287.038 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 59.2579 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 289.419 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.5608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.128 LAYER met4  ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 61.7425 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 302.807 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.981399 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.5000 0.4850 156.6400 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 62.3286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 333.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 66.0549 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 339.4 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 153.4400 0.4850 153.5800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.5035 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 302.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 66.4023 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 315.943 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.756604 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 150.3800 0.4850 150.5200 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.0154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 46.3239 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 210.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.898113 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.3200 0.4850 147.4600 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.2031 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 60.534 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 279.35 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.630818 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 144.2600 0.4850 144.4000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.9 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 282.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.6828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 30.9923 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 97.4731 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.60386 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 141.2000 0.4850 141.3400 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.9606 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 32.9482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 164.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.463989 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.1400 0.4850 138.2800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0655 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met2  ;
    ANTENNAMAXAREACAR 44.0147 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 209.6 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.672557 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.1635 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.128 LAYER met3  ;
    ANTENNAGATEAREA 2.6505 LAYER met3  ;
    ANTENNAMAXAREACAR 52.3767 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 254.546 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.687649 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.7356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.864 LAYER met4  ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 60.4265 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.751 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.687649 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.0800 0.4850 135.2200 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met2  ;
    ANTENNAMAXAREACAR 25.0722 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.361 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.484591 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.9298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.896 LAYER met3  ;
    ANTENNAGATEAREA 1.908 LAYER met3  ;
    ANTENNAMAXAREACAR 50.2779 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 239.166 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.597874 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.6486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.4 LAYER met4  ;
    ANTENNAGATEAREA 3.6045 LAYER met4  ;
    ANTENNAMAXAREACAR 57.1162 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 275.898 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.598421 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 56.6089 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.621 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.60386 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.9600 0.4850 129.1000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 55.3128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 295.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 48.2364 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 241.987 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.9000 0.4850 126.0400 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.292 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met2  ;
    ANTENNAMAXAREACAR 41.3327 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 194.469 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.544744 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.6714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.512 LAYER met3  ;
    ANTENNAGATEAREA 3.4455 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3638 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 237.572 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 122.8400 0.4850 122.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5625 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.4038 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.906 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 23.9195 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.258 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9481 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.6 LAYER met4  ;
    ANTENNAGATEAREA 3.6045 LAYER met4  ;
    ANTENNAMAXAREACAR 52.4094 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.504 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.1675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 195.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.6608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.328 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 214.3000 230.4600 214.4400 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.272 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 211.5800 230.4600 211.7200 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.0798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 304.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 208.5200 230.4600 208.6600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.293 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.2258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 205.4600 230.4600 205.6000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.3308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 202.4000 230.4600 202.5400 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.4578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 199.3400 230.4600 199.4800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.7566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.976 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 196.2800 230.4600 196.4200 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 193.2200 230.4600 193.3600 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.7248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 340.336 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 190.1600 230.4600 190.3000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.077 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 187.1000 230.4600 187.2400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.3952 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 184.0400 230.4600 184.1800 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.6128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.7766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 180.9800 230.4600 181.1200 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.055 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 177.9200 230.4600 178.0600 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.462 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.7024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 174.8600 230.4600 175.0000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.1194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.048 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 171.8000 230.4600 171.9400 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.4062 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.048 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 168.7400 230.4600 168.8800 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 165.6800 230.4600 165.8200 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.42 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 162.6200 230.4600 162.7600 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.1836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.92 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 159.5600 230.4600 159.7000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.9498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 156.5000 230.4600 156.6400 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 153.4400 230.4600 153.5800 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 150.3800 230.4600 150.5200 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.81 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 147.3200 230.4600 147.4600 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.353 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.7538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 144.2600 230.4600 144.4000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.586 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 141.2000 230.4600 141.3400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.89 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 138.1400 230.4600 138.2800 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 244.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 135.0800 230.4600 135.2200 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 132.0200 230.4600 132.1600 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 128.9600 230.4600 129.1000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.072 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 125.9000 230.4600 126.0400 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.312 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 263.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.1398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 122.8400 230.4600 122.9800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 120.1200 230.4600 120.2600 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.9995 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3832 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.4997 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.112097 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 214.0600 0.0000 214.2000 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.723 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.5798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 24.0181 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 90.3538 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.399033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.4600 0.0000 209.6000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.886 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.6418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 238.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met3  ;
    ANTENNAMAXAREACAR 31.7739 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.398 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.446448 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 204.4000 0.0000 204.5400 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.91 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.3618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 39.0787 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.033 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.461539 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 199.3400 0.0000 199.4800 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.1788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 30.5002 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.24 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.454309 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 193.8200 0.0000 193.9600 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.572 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.3246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met3  ;
    ANTENNAMAXAREACAR 64.9955 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 318.061 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.496226 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 189.6800 0.0000 189.8200 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.358 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5771 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.4716 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.405716 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8442 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.1276 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.425572 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 17.9848 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 68.5534 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.425572 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 184.6200 0.0000 184.7600 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.7115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met2  ;
    ANTENNAMAXAREACAR 13.6523 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.0659 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.272372 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.7768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.28 LAYER met3  ;
    ANTENNAGATEAREA 3.2865 LAYER met3  ;
    ANTENNAMAXAREACAR 15.41 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 53.5836 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354717 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 179.5600 0.0000 179.7000 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8516 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.954 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.4641 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.281533 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.9607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.256 LAYER met3  ;
    ANTENNAGATEAREA 3.2865 LAYER met3  ;
    ANTENNAMAXAREACAR 17.4847 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.5829 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.386164 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 174.5000 0.0000 174.6400 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.9028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 45.1894 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.552 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.502108 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.4400 0.0000 169.5800 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.0695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7093 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.8973 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.389251 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 164.8400 0.0000 164.9800 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.574 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.9296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 47.7566 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.974 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.544204 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 159.7800 0.0000 159.9200 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 19.138 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 80.5785 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.493996 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 154.7200 0.0000 154.8600 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.804 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.4584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 27.946 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 92.4916 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.529373 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 149.6600 0.0000 149.8000 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.8698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 32.4788 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 140.828 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.644931 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 144.1400 0.0000 144.2800 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.4818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6611 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 98.1096 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.472464 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 140.0000 0.0000 140.1400 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.081 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.0828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 72.0867 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 141.763 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.577065 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 134.9400 0.0000 135.0800 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.9966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2044 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 143.599 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.494667 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 129.4200 0.0000 129.5600 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.2898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 40.5596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.559062 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 124.8200 0.0000 124.9600 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.2314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 34.8935 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 157.987 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.730398 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 120.2200 0.0000 120.3600 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.48 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.239 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.6108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 214.0600 229.3550 214.2000 229.8400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.129 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 205.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.9918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.76 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.4600 229.3550 209.6000 229.8400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.2866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.136 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 204.4000 229.3550 204.5400 229.8400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.3400 229.3550 199.4800 229.8400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.96 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 194.2800 229.3550 194.4200 229.8400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.3738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 189.6800 229.3550 189.8200 229.8400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.867 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.7638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.544 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 184.6200 229.3550 184.7600 229.8400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.032 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.5308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 179.5600 229.3550 179.7000 229.8400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.696 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.2978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 174.5000 229.3550 174.6400 229.8400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.7318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 169.4400 229.3550 169.5800 229.8400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.6158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 345.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.8400 229.3550 164.9800 229.8400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.532 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 159.7800 229.3550 159.9200 229.8400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 154.7200 229.3550 154.8600 229.8400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.676 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.3386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 149.2000 229.3550 149.3400 229.8400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.867 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.1108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 144.6000 229.3550 144.7400 229.8400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.3768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 139.5400 229.3550 139.6800 229.8400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.4800 229.3550 134.6200 229.8400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.8800 229.3550 130.0200 229.8400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7747 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.8200 229.3550 124.9600 229.8400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.7155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.2200 229.3550 120.3600 229.8400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 190.1200 5.4300 191.7200 224.0700 ;
        RECT 160.1200 5.4300 161.7200 224.0700 ;
        RECT 130.1200 5.4300 131.7200 224.0700 ;
        RECT 100.1200 5.4300 101.7200 224.0700 ;
        RECT 70.1200 5.4300 71.7200 224.0700 ;
        RECT 40.1200 5.4300 41.7200 224.0700 ;
        RECT 221.9000 5.4300 224.9000 224.0700 ;
        RECT 5.5600 5.4300 8.5600 224.0700 ;
      LAYER met3 ;
        RECT 5.5600 5.4300 224.9000 8.4300 ;
        RECT 5.5600 221.0700 224.9000 224.0700 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 193.3200 1.4300 194.9200 228.0700 ;
        RECT 163.3200 1.4300 164.9200 228.0700 ;
        RECT 133.3200 1.4300 134.9200 228.0700 ;
        RECT 103.3200 1.4300 104.9200 228.0700 ;
        RECT 73.3200 1.4300 74.9200 228.0700 ;
        RECT 43.3200 1.4300 44.9200 228.0700 ;
        RECT 13.3200 1.4300 14.9200 228.0700 ;
        RECT 225.9000 1.4300 228.9000 228.0700 ;
        RECT 1.5600 1.4300 4.5600 228.0700 ;
      LAYER met3 ;
        RECT 1.5600 1.4300 228.9000 4.4300 ;
        RECT 1.5600 225.0700 228.9000 228.0700 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 109.9650 229.3400 230.4600 229.8400 ;
      RECT 108.5850 229.3400 109.4550 229.8400 ;
      RECT 107.2050 229.3400 108.0750 229.8400 ;
      RECT 105.8250 229.3400 106.6950 229.8400 ;
      RECT 104.4450 229.3400 105.3150 229.8400 ;
      RECT 103.0650 229.3400 103.9350 229.8400 ;
      RECT 101.6850 229.3400 102.5550 229.8400 ;
      RECT 100.3050 229.3400 101.1750 229.8400 ;
      RECT 98.9250 229.3400 99.7950 229.8400 ;
      RECT 98.0050 229.3400 98.4150 229.8400 ;
      RECT 96.6250 229.3400 97.4950 229.8400 ;
      RECT 95.2450 229.3400 96.1150 229.8400 ;
      RECT 93.8650 229.3400 94.7350 229.8400 ;
      RECT 92.4850 229.3400 93.3550 229.8400 ;
      RECT 91.1050 229.3400 91.9750 229.8400 ;
      RECT 89.7250 229.3400 90.5950 229.8400 ;
      RECT 88.3450 229.3400 89.2150 229.8400 ;
      RECT 86.9650 229.3400 87.8350 229.8400 ;
      RECT 86.0450 229.3400 86.4550 229.8400 ;
      RECT 84.6650 229.3400 85.5350 229.8400 ;
      RECT 83.2850 229.3400 84.1550 229.8400 ;
      RECT 81.9050 229.3400 82.7750 229.8400 ;
      RECT 80.5250 229.3400 81.3950 229.8400 ;
      RECT 79.1450 229.3400 80.0150 229.8400 ;
      RECT 77.7650 229.3400 78.6350 229.8400 ;
      RECT 76.3850 229.3400 77.2550 229.8400 ;
      RECT 75.0050 229.3400 75.8750 229.8400 ;
      RECT 74.0850 229.3400 74.4950 229.8400 ;
      RECT 72.7050 229.3400 73.5750 229.8400 ;
      RECT 71.3250 229.3400 72.1950 229.8400 ;
      RECT 69.9450 229.3400 70.8150 229.8400 ;
      RECT 68.5650 229.3400 69.4350 229.8400 ;
      RECT 67.1850 229.3400 68.0550 229.8400 ;
      RECT 65.8050 229.3400 66.6750 229.8400 ;
      RECT 64.4250 229.3400 65.2950 229.8400 ;
      RECT 63.0450 229.3400 63.9150 229.8400 ;
      RECT 62.1250 229.3400 62.5350 229.8400 ;
      RECT 60.7450 229.3400 61.6150 229.8400 ;
      RECT 59.3650 229.3400 60.2350 229.8400 ;
      RECT 57.9850 229.3400 58.8550 229.8400 ;
      RECT 56.6050 229.3400 57.4750 229.8400 ;
      RECT 55.2250 229.3400 56.0950 229.8400 ;
      RECT 53.8450 229.3400 54.7150 229.8400 ;
      RECT 52.4650 229.3400 53.3350 229.8400 ;
      RECT 51.0850 229.3400 51.9550 229.8400 ;
      RECT 50.1650 229.3400 50.5750 229.8400 ;
      RECT 48.7850 229.3400 49.6550 229.8400 ;
      RECT 47.4050 229.3400 48.2750 229.8400 ;
      RECT 46.0250 229.3400 46.8950 229.8400 ;
      RECT 44.6450 229.3400 45.5150 229.8400 ;
      RECT 43.2650 229.3400 44.1350 229.8400 ;
      RECT 41.8850 229.3400 42.7550 229.8400 ;
      RECT 40.5050 229.3400 41.3750 229.8400 ;
      RECT 39.1250 229.3400 39.9950 229.8400 ;
      RECT 38.2050 229.3400 38.6150 229.8400 ;
      RECT 36.8250 229.3400 37.6950 229.8400 ;
      RECT 35.4450 229.3400 36.3150 229.8400 ;
      RECT 34.0650 229.3400 34.9350 229.8400 ;
      RECT 32.6850 229.3400 33.5550 229.8400 ;
      RECT 31.3050 229.3400 32.1750 229.8400 ;
      RECT 29.9250 229.3400 30.7950 229.8400 ;
      RECT 28.5450 229.3400 29.4150 229.8400 ;
      RECT 27.1650 229.3400 28.0350 229.8400 ;
      RECT 26.2450 229.3400 26.6550 229.8400 ;
      RECT 24.8650 229.3400 25.7350 229.8400 ;
      RECT 23.4850 229.3400 24.3550 229.8400 ;
      RECT 22.1050 229.3400 22.9750 229.8400 ;
      RECT 20.7250 229.3400 21.5950 229.8400 ;
      RECT 19.3450 229.3400 20.2150 229.8400 ;
      RECT 17.9650 229.3400 18.8350 229.8400 ;
      RECT 16.5850 229.3400 17.4550 229.8400 ;
      RECT 15.6650 229.3400 16.0750 229.8400 ;
      RECT 0.0000 229.3400 15.1550 229.8400 ;
      RECT 0.0000 0.5000 230.4600 229.3400 ;
      RECT 109.9650 0.0000 230.4600 0.5000 ;
      RECT 108.5850 0.0000 109.4550 0.5000 ;
      RECT 107.2050 0.0000 108.0750 0.5000 ;
      RECT 105.8250 0.0000 106.6950 0.5000 ;
      RECT 104.4450 0.0000 105.3150 0.5000 ;
      RECT 103.0650 0.0000 103.9350 0.5000 ;
      RECT 101.6850 0.0000 102.5550 0.5000 ;
      RECT 100.3050 0.0000 101.1750 0.5000 ;
      RECT 98.9250 0.0000 99.7950 0.5000 ;
      RECT 98.0050 0.0000 98.4150 0.5000 ;
      RECT 96.6250 0.0000 97.4950 0.5000 ;
      RECT 95.2450 0.0000 96.1150 0.5000 ;
      RECT 93.8650 0.0000 94.7350 0.5000 ;
      RECT 92.4850 0.0000 93.3550 0.5000 ;
      RECT 91.1050 0.0000 91.9750 0.5000 ;
      RECT 89.7250 0.0000 90.5950 0.5000 ;
      RECT 88.3450 0.0000 89.2150 0.5000 ;
      RECT 86.9650 0.0000 87.8350 0.5000 ;
      RECT 86.0450 0.0000 86.4550 0.5000 ;
      RECT 84.6650 0.0000 85.5350 0.5000 ;
      RECT 83.2850 0.0000 84.1550 0.5000 ;
      RECT 81.9050 0.0000 82.7750 0.5000 ;
      RECT 80.5250 0.0000 81.3950 0.5000 ;
      RECT 79.1450 0.0000 80.0150 0.5000 ;
      RECT 77.7650 0.0000 78.6350 0.5000 ;
      RECT 76.3850 0.0000 77.2550 0.5000 ;
      RECT 75.0050 0.0000 75.8750 0.5000 ;
      RECT 74.0850 0.0000 74.4950 0.5000 ;
      RECT 72.7050 0.0000 73.5750 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 69.9450 0.0000 70.8150 0.5000 ;
      RECT 68.5650 0.0000 69.4350 0.5000 ;
      RECT 67.1850 0.0000 68.0550 0.5000 ;
      RECT 65.8050 0.0000 66.6750 0.5000 ;
      RECT 64.4250 0.0000 65.2950 0.5000 ;
      RECT 63.0450 0.0000 63.9150 0.5000 ;
      RECT 62.1250 0.0000 62.5350 0.5000 ;
      RECT 60.7450 0.0000 61.6150 0.5000 ;
      RECT 59.3650 0.0000 60.2350 0.5000 ;
      RECT 57.9850 0.0000 58.8550 0.5000 ;
      RECT 56.6050 0.0000 57.4750 0.5000 ;
      RECT 55.2250 0.0000 56.0950 0.5000 ;
      RECT 53.8450 0.0000 54.7150 0.5000 ;
      RECT 52.4650 0.0000 53.3350 0.5000 ;
      RECT 51.0850 0.0000 51.9550 0.5000 ;
      RECT 50.1650 0.0000 50.5750 0.5000 ;
      RECT 48.7850 0.0000 49.6550 0.5000 ;
      RECT 47.4050 0.0000 48.2750 0.5000 ;
      RECT 46.0250 0.0000 46.8950 0.5000 ;
      RECT 44.6450 0.0000 45.5150 0.5000 ;
      RECT 43.2650 0.0000 44.1350 0.5000 ;
      RECT 41.8850 0.0000 42.7550 0.5000 ;
      RECT 40.5050 0.0000 41.3750 0.5000 ;
      RECT 39.1250 0.0000 39.9950 0.5000 ;
      RECT 38.2050 0.0000 38.6150 0.5000 ;
      RECT 36.8250 0.0000 37.6950 0.5000 ;
      RECT 35.4450 0.0000 36.3150 0.5000 ;
      RECT 34.0650 0.0000 34.9350 0.5000 ;
      RECT 32.6850 0.0000 33.5550 0.5000 ;
      RECT 31.3050 0.0000 32.1750 0.5000 ;
      RECT 29.9250 0.0000 30.7950 0.5000 ;
      RECT 28.5450 0.0000 29.4150 0.5000 ;
      RECT 27.1650 0.0000 28.0350 0.5000 ;
      RECT 26.2450 0.0000 26.6550 0.5000 ;
      RECT 24.8650 0.0000 25.7350 0.5000 ;
      RECT 23.4850 0.0000 24.3550 0.5000 ;
      RECT 22.1050 0.0000 22.9750 0.5000 ;
      RECT 20.7250 0.0000 21.5950 0.5000 ;
      RECT 19.3450 0.0000 20.2150 0.5000 ;
      RECT 17.9650 0.0000 18.8350 0.5000 ;
      RECT 16.5850 0.0000 17.4550 0.5000 ;
      RECT 15.6650 0.0000 16.0750 0.5000 ;
      RECT 0.0000 0.0000 15.1550 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 230.4600 229.8400 ;
    LAYER met2 ;
      RECT 214.3400 229.2150 230.4600 229.8400 ;
      RECT 209.7400 229.2150 213.9200 229.8400 ;
      RECT 204.6800 229.2150 209.3200 229.8400 ;
      RECT 199.6200 229.2150 204.2600 229.8400 ;
      RECT 194.5600 229.2150 199.2000 229.8400 ;
      RECT 189.9600 229.2150 194.1400 229.8400 ;
      RECT 184.9000 229.2150 189.5400 229.8400 ;
      RECT 179.8400 229.2150 184.4800 229.8400 ;
      RECT 174.7800 229.2150 179.4200 229.8400 ;
      RECT 169.7200 229.2150 174.3600 229.8400 ;
      RECT 165.1200 229.2150 169.3000 229.8400 ;
      RECT 160.0600 229.2150 164.7000 229.8400 ;
      RECT 155.0000 229.2150 159.6400 229.8400 ;
      RECT 149.4800 229.2150 154.5800 229.8400 ;
      RECT 144.8800 229.2150 149.0600 229.8400 ;
      RECT 139.8200 229.2150 144.4600 229.8400 ;
      RECT 134.7600 229.2150 139.4000 229.8400 ;
      RECT 130.1600 229.2150 134.3400 229.8400 ;
      RECT 125.1000 229.2150 129.7400 229.8400 ;
      RECT 120.5000 229.2150 124.6800 229.8400 ;
      RECT 0.0000 229.2150 120.0800 229.8400 ;
      RECT 0.0000 228.2100 230.4600 229.2150 ;
      RECT 195.0600 224.2100 225.7600 228.2100 ;
      RECT 165.0600 224.2100 193.1800 228.2100 ;
      RECT 135.0600 224.2100 163.1800 228.2100 ;
      RECT 105.0600 224.2100 133.1800 228.2100 ;
      RECT 75.0600 224.2100 103.1800 228.2100 ;
      RECT 45.0600 224.2100 73.1800 228.2100 ;
      RECT 15.0600 224.2100 43.1800 228.2100 ;
      RECT 4.7000 224.2100 13.1800 228.2100 ;
      RECT 229.0400 214.5800 230.4600 228.2100 ;
      RECT 0.0000 214.5800 1.4200 228.2100 ;
      RECT 229.0400 214.1600 229.8350 214.5800 ;
      RECT 0.6250 214.1600 1.4200 214.5800 ;
      RECT 229.0400 211.8600 230.4600 214.1600 ;
      RECT 0.0000 211.8600 1.4200 214.1600 ;
      RECT 229.0400 211.4400 229.8350 211.8600 ;
      RECT 0.6250 211.4400 1.4200 211.8600 ;
      RECT 229.0400 208.8000 230.4600 211.4400 ;
      RECT 0.0000 208.8000 1.4200 211.4400 ;
      RECT 229.0400 208.3800 229.8350 208.8000 ;
      RECT 0.6250 208.3800 1.4200 208.8000 ;
      RECT 229.0400 205.7400 230.4600 208.3800 ;
      RECT 0.0000 205.7400 1.4200 208.3800 ;
      RECT 229.0400 205.3200 229.8350 205.7400 ;
      RECT 0.6250 205.3200 1.4200 205.7400 ;
      RECT 229.0400 202.6800 230.4600 205.3200 ;
      RECT 0.0000 202.6800 1.4200 205.3200 ;
      RECT 229.0400 202.2600 229.8350 202.6800 ;
      RECT 0.6250 202.2600 1.4200 202.6800 ;
      RECT 229.0400 199.6200 230.4600 202.2600 ;
      RECT 0.0000 199.6200 1.4200 202.2600 ;
      RECT 229.0400 199.2000 229.8350 199.6200 ;
      RECT 0.6250 199.2000 1.4200 199.6200 ;
      RECT 229.0400 196.5600 230.4600 199.2000 ;
      RECT 0.0000 196.5600 1.4200 199.2000 ;
      RECT 229.0400 196.1400 229.8350 196.5600 ;
      RECT 0.6250 196.1400 1.4200 196.5600 ;
      RECT 229.0400 193.5000 230.4600 196.1400 ;
      RECT 0.0000 193.5000 1.4200 196.1400 ;
      RECT 229.0400 193.0800 229.8350 193.5000 ;
      RECT 0.6250 193.0800 1.4200 193.5000 ;
      RECT 229.0400 190.4400 230.4600 193.0800 ;
      RECT 0.0000 190.4400 1.4200 193.0800 ;
      RECT 229.0400 190.0200 229.8350 190.4400 ;
      RECT 0.6250 190.0200 1.4200 190.4400 ;
      RECT 229.0400 187.3800 230.4600 190.0200 ;
      RECT 0.0000 187.3800 1.4200 190.0200 ;
      RECT 229.0400 186.9600 229.8350 187.3800 ;
      RECT 0.6250 186.9600 1.4200 187.3800 ;
      RECT 229.0400 184.3200 230.4600 186.9600 ;
      RECT 0.0000 184.3200 1.4200 186.9600 ;
      RECT 229.0400 183.9000 229.8350 184.3200 ;
      RECT 0.6250 183.9000 1.4200 184.3200 ;
      RECT 229.0400 181.2600 230.4600 183.9000 ;
      RECT 0.0000 181.2600 1.4200 183.9000 ;
      RECT 229.0400 180.8400 229.8350 181.2600 ;
      RECT 0.6250 180.8400 1.4200 181.2600 ;
      RECT 229.0400 178.2000 230.4600 180.8400 ;
      RECT 0.0000 178.2000 1.4200 180.8400 ;
      RECT 229.0400 177.7800 229.8350 178.2000 ;
      RECT 0.6250 177.7800 1.4200 178.2000 ;
      RECT 229.0400 175.1400 230.4600 177.7800 ;
      RECT 0.0000 175.1400 1.4200 177.7800 ;
      RECT 229.0400 174.7200 229.8350 175.1400 ;
      RECT 0.6250 174.7200 1.4200 175.1400 ;
      RECT 229.0400 172.0800 230.4600 174.7200 ;
      RECT 0.0000 172.0800 1.4200 174.7200 ;
      RECT 229.0400 171.6600 229.8350 172.0800 ;
      RECT 0.6250 171.6600 1.4200 172.0800 ;
      RECT 229.0400 169.0200 230.4600 171.6600 ;
      RECT 0.0000 169.0200 1.4200 171.6600 ;
      RECT 229.0400 168.6000 229.8350 169.0200 ;
      RECT 0.6250 168.6000 1.4200 169.0200 ;
      RECT 229.0400 165.9600 230.4600 168.6000 ;
      RECT 0.0000 165.9600 1.4200 168.6000 ;
      RECT 229.0400 165.5400 229.8350 165.9600 ;
      RECT 0.6250 165.5400 1.4200 165.9600 ;
      RECT 229.0400 162.9000 230.4600 165.5400 ;
      RECT 0.0000 162.9000 1.4200 165.5400 ;
      RECT 229.0400 162.4800 229.8350 162.9000 ;
      RECT 0.6250 162.4800 1.4200 162.9000 ;
      RECT 229.0400 159.8400 230.4600 162.4800 ;
      RECT 0.0000 159.8400 1.4200 162.4800 ;
      RECT 229.0400 159.4200 229.8350 159.8400 ;
      RECT 0.6250 159.4200 1.4200 159.8400 ;
      RECT 229.0400 156.7800 230.4600 159.4200 ;
      RECT 0.0000 156.7800 1.4200 159.4200 ;
      RECT 229.0400 156.3600 229.8350 156.7800 ;
      RECT 0.6250 156.3600 1.4200 156.7800 ;
      RECT 229.0400 153.7200 230.4600 156.3600 ;
      RECT 0.0000 153.7200 1.4200 156.3600 ;
      RECT 229.0400 153.3000 229.8350 153.7200 ;
      RECT 0.6250 153.3000 1.4200 153.7200 ;
      RECT 229.0400 150.6600 230.4600 153.3000 ;
      RECT 0.0000 150.6600 1.4200 153.3000 ;
      RECT 229.0400 150.2400 229.8350 150.6600 ;
      RECT 0.6250 150.2400 1.4200 150.6600 ;
      RECT 229.0400 147.6000 230.4600 150.2400 ;
      RECT 0.0000 147.6000 1.4200 150.2400 ;
      RECT 229.0400 147.1800 229.8350 147.6000 ;
      RECT 0.6250 147.1800 1.4200 147.6000 ;
      RECT 229.0400 144.5400 230.4600 147.1800 ;
      RECT 0.0000 144.5400 1.4200 147.1800 ;
      RECT 229.0400 144.1200 229.8350 144.5400 ;
      RECT 0.6250 144.1200 1.4200 144.5400 ;
      RECT 229.0400 141.4800 230.4600 144.1200 ;
      RECT 0.0000 141.4800 1.4200 144.1200 ;
      RECT 229.0400 141.0600 229.8350 141.4800 ;
      RECT 0.6250 141.0600 1.4200 141.4800 ;
      RECT 229.0400 138.4200 230.4600 141.0600 ;
      RECT 0.0000 138.4200 1.4200 141.0600 ;
      RECT 229.0400 138.0000 229.8350 138.4200 ;
      RECT 0.6250 138.0000 1.4200 138.4200 ;
      RECT 229.0400 135.3600 230.4600 138.0000 ;
      RECT 0.0000 135.3600 1.4200 138.0000 ;
      RECT 229.0400 134.9400 229.8350 135.3600 ;
      RECT 0.6250 134.9400 1.4200 135.3600 ;
      RECT 229.0400 132.3000 230.4600 134.9400 ;
      RECT 0.0000 132.3000 1.4200 134.9400 ;
      RECT 229.0400 131.8800 229.8350 132.3000 ;
      RECT 0.6250 131.8800 1.4200 132.3000 ;
      RECT 229.0400 129.2400 230.4600 131.8800 ;
      RECT 0.0000 129.2400 1.4200 131.8800 ;
      RECT 229.0400 128.8200 229.8350 129.2400 ;
      RECT 0.6250 128.8200 1.4200 129.2400 ;
      RECT 229.0400 126.1800 230.4600 128.8200 ;
      RECT 0.0000 126.1800 1.4200 128.8200 ;
      RECT 229.0400 125.7600 229.8350 126.1800 ;
      RECT 0.6250 125.7600 1.4200 126.1800 ;
      RECT 229.0400 123.1200 230.4600 125.7600 ;
      RECT 0.0000 123.1200 1.4200 125.7600 ;
      RECT 229.0400 122.7000 229.8350 123.1200 ;
      RECT 0.6250 122.7000 1.4200 123.1200 ;
      RECT 229.0400 120.4000 230.4600 122.7000 ;
      RECT 0.0000 120.4000 1.4200 122.7000 ;
      RECT 229.0400 119.9800 229.8350 120.4000 ;
      RECT 0.6250 119.9800 1.4200 120.4000 ;
      RECT 229.0400 109.8600 230.4600 119.9800 ;
      RECT 0.0000 109.8600 1.4200 119.9800 ;
      RECT 229.0400 109.4400 229.8350 109.8600 ;
      RECT 0.6250 109.4400 1.4200 109.8600 ;
      RECT 229.0400 108.5000 230.4600 109.4400 ;
      RECT 0.0000 108.5000 1.4200 109.4400 ;
      RECT 229.0400 108.0800 229.8350 108.5000 ;
      RECT 0.6250 108.0800 1.4200 108.5000 ;
      RECT 229.0400 107.1400 230.4600 108.0800 ;
      RECT 0.0000 107.1400 1.4200 108.0800 ;
      RECT 229.0400 106.7200 229.8350 107.1400 ;
      RECT 0.6250 106.7200 1.4200 107.1400 ;
      RECT 229.0400 105.4400 230.4600 106.7200 ;
      RECT 0.0000 105.4400 1.4200 106.7200 ;
      RECT 229.0400 105.0200 229.8350 105.4400 ;
      RECT 0.6250 105.0200 1.4200 105.4400 ;
      RECT 229.0400 104.0800 230.4600 105.0200 ;
      RECT 0.0000 104.0800 1.4200 105.0200 ;
      RECT 229.0400 103.6600 229.8350 104.0800 ;
      RECT 0.6250 103.6600 1.4200 104.0800 ;
      RECT 229.0400 102.3800 230.4600 103.6600 ;
      RECT 0.0000 102.3800 1.4200 103.6600 ;
      RECT 229.0400 101.9600 229.8350 102.3800 ;
      RECT 0.6250 101.9600 1.4200 102.3800 ;
      RECT 229.0400 101.0200 230.4600 101.9600 ;
      RECT 0.0000 101.0200 1.4200 101.9600 ;
      RECT 229.0400 100.6000 229.8350 101.0200 ;
      RECT 0.6250 100.6000 1.4200 101.0200 ;
      RECT 229.0400 99.3200 230.4600 100.6000 ;
      RECT 0.0000 99.3200 1.4200 100.6000 ;
      RECT 229.0400 98.9000 229.8350 99.3200 ;
      RECT 0.6250 98.9000 1.4200 99.3200 ;
      RECT 229.0400 97.9600 230.4600 98.9000 ;
      RECT 0.0000 97.9600 1.4200 98.9000 ;
      RECT 229.0400 97.5400 229.8350 97.9600 ;
      RECT 0.6250 97.5400 1.4200 97.9600 ;
      RECT 229.0400 96.6000 230.4600 97.5400 ;
      RECT 0.0000 96.6000 1.4200 97.5400 ;
      RECT 229.0400 96.1800 229.8350 96.6000 ;
      RECT 0.6250 96.1800 1.4200 96.6000 ;
      RECT 229.0400 94.9000 230.4600 96.1800 ;
      RECT 0.0000 94.9000 1.4200 96.1800 ;
      RECT 229.0400 94.4800 229.8350 94.9000 ;
      RECT 0.6250 94.4800 1.4200 94.9000 ;
      RECT 229.0400 93.5400 230.4600 94.4800 ;
      RECT 0.0000 93.5400 1.4200 94.4800 ;
      RECT 229.0400 93.1200 229.8350 93.5400 ;
      RECT 0.6250 93.1200 1.4200 93.5400 ;
      RECT 229.0400 91.8400 230.4600 93.1200 ;
      RECT 0.0000 91.8400 1.4200 93.1200 ;
      RECT 229.0400 91.4200 229.8350 91.8400 ;
      RECT 0.6250 91.4200 1.4200 91.8400 ;
      RECT 229.0400 90.4800 230.4600 91.4200 ;
      RECT 0.0000 90.4800 1.4200 91.4200 ;
      RECT 229.0400 90.0600 229.8350 90.4800 ;
      RECT 0.6250 90.0600 1.4200 90.4800 ;
      RECT 229.0400 88.7800 230.4600 90.0600 ;
      RECT 0.0000 88.7800 1.4200 90.0600 ;
      RECT 229.0400 88.3600 229.8350 88.7800 ;
      RECT 0.6250 88.3600 1.4200 88.7800 ;
      RECT 229.0400 87.4200 230.4600 88.3600 ;
      RECT 0.0000 87.4200 1.4200 88.3600 ;
      RECT 229.0400 87.0000 229.8350 87.4200 ;
      RECT 0.6250 87.0000 1.4200 87.4200 ;
      RECT 229.0400 86.0600 230.4600 87.0000 ;
      RECT 0.0000 86.0600 1.4200 87.0000 ;
      RECT 229.0400 85.6400 229.8350 86.0600 ;
      RECT 0.6250 85.6400 1.4200 86.0600 ;
      RECT 229.0400 84.3600 230.4600 85.6400 ;
      RECT 0.0000 84.3600 1.4200 85.6400 ;
      RECT 229.0400 83.9400 229.8350 84.3600 ;
      RECT 0.6250 83.9400 1.4200 84.3600 ;
      RECT 229.0400 83.0000 230.4600 83.9400 ;
      RECT 0.0000 83.0000 1.4200 83.9400 ;
      RECT 229.0400 82.5800 229.8350 83.0000 ;
      RECT 0.6250 82.5800 1.4200 83.0000 ;
      RECT 229.0400 81.3000 230.4600 82.5800 ;
      RECT 0.0000 81.3000 1.4200 82.5800 ;
      RECT 229.0400 80.8800 229.8350 81.3000 ;
      RECT 0.6250 80.8800 1.4200 81.3000 ;
      RECT 229.0400 79.9400 230.4600 80.8800 ;
      RECT 0.0000 79.9400 1.4200 80.8800 ;
      RECT 229.0400 79.5200 229.8350 79.9400 ;
      RECT 0.6250 79.5200 1.4200 79.9400 ;
      RECT 229.0400 78.2400 230.4600 79.5200 ;
      RECT 0.0000 78.2400 1.4200 79.5200 ;
      RECT 229.0400 77.8200 229.8350 78.2400 ;
      RECT 0.6250 77.8200 1.4200 78.2400 ;
      RECT 229.0400 76.8800 230.4600 77.8200 ;
      RECT 0.0000 76.8800 1.4200 77.8200 ;
      RECT 229.0400 76.4600 229.8350 76.8800 ;
      RECT 0.6250 76.4600 1.4200 76.8800 ;
      RECT 229.0400 75.5200 230.4600 76.4600 ;
      RECT 0.0000 75.5200 1.4200 76.4600 ;
      RECT 229.0400 75.1000 229.8350 75.5200 ;
      RECT 0.6250 75.1000 1.4200 75.5200 ;
      RECT 229.0400 73.8200 230.4600 75.1000 ;
      RECT 0.0000 73.8200 1.4200 75.1000 ;
      RECT 229.0400 73.4000 229.8350 73.8200 ;
      RECT 0.6250 73.4000 1.4200 73.8200 ;
      RECT 229.0400 72.4600 230.4600 73.4000 ;
      RECT 0.0000 72.4600 1.4200 73.4000 ;
      RECT 229.0400 72.0400 229.8350 72.4600 ;
      RECT 0.6250 72.0400 1.4200 72.4600 ;
      RECT 229.0400 70.7600 230.4600 72.0400 ;
      RECT 0.0000 70.7600 1.4200 72.0400 ;
      RECT 229.0400 70.3400 229.8350 70.7600 ;
      RECT 0.6250 70.3400 1.4200 70.7600 ;
      RECT 229.0400 69.4000 230.4600 70.3400 ;
      RECT 0.0000 69.4000 1.4200 70.3400 ;
      RECT 229.0400 68.9800 229.8350 69.4000 ;
      RECT 0.6250 68.9800 1.4200 69.4000 ;
      RECT 229.0400 67.7000 230.4600 68.9800 ;
      RECT 0.0000 67.7000 1.4200 68.9800 ;
      RECT 229.0400 67.2800 229.8350 67.7000 ;
      RECT 0.6250 67.2800 1.4200 67.7000 ;
      RECT 229.0400 66.3400 230.4600 67.2800 ;
      RECT 0.0000 66.3400 1.4200 67.2800 ;
      RECT 229.0400 65.9200 229.8350 66.3400 ;
      RECT 0.6250 65.9200 1.4200 66.3400 ;
      RECT 229.0400 64.9800 230.4600 65.9200 ;
      RECT 0.0000 64.9800 1.4200 65.9200 ;
      RECT 229.0400 64.5600 229.8350 64.9800 ;
      RECT 0.6250 64.5600 1.4200 64.9800 ;
      RECT 229.0400 63.2800 230.4600 64.5600 ;
      RECT 0.0000 63.2800 1.4200 64.5600 ;
      RECT 229.0400 62.8600 229.8350 63.2800 ;
      RECT 0.6250 62.8600 1.4200 63.2800 ;
      RECT 229.0400 61.9200 230.4600 62.8600 ;
      RECT 0.0000 61.9200 1.4200 62.8600 ;
      RECT 229.0400 61.5000 229.8350 61.9200 ;
      RECT 0.6250 61.5000 1.4200 61.9200 ;
      RECT 229.0400 60.2200 230.4600 61.5000 ;
      RECT 0.0000 60.2200 1.4200 61.5000 ;
      RECT 229.0400 59.8000 229.8350 60.2200 ;
      RECT 0.6250 59.8000 1.4200 60.2200 ;
      RECT 229.0400 58.8600 230.4600 59.8000 ;
      RECT 0.0000 58.8600 1.4200 59.8000 ;
      RECT 229.0400 58.4400 229.8350 58.8600 ;
      RECT 0.6250 58.4400 1.4200 58.8600 ;
      RECT 229.0400 57.5000 230.4600 58.4400 ;
      RECT 0.0000 57.5000 1.4200 58.4400 ;
      RECT 229.0400 57.0800 229.8350 57.5000 ;
      RECT 0.6250 57.0800 1.4200 57.5000 ;
      RECT 229.0400 55.8000 230.4600 57.0800 ;
      RECT 0.0000 55.8000 1.4200 57.0800 ;
      RECT 229.0400 55.3800 229.8350 55.8000 ;
      RECT 0.6250 55.3800 1.4200 55.8000 ;
      RECT 229.0400 54.4400 230.4600 55.3800 ;
      RECT 0.0000 54.4400 1.4200 55.3800 ;
      RECT 229.0400 54.0200 229.8350 54.4400 ;
      RECT 0.6250 54.0200 1.4200 54.4400 ;
      RECT 229.0400 52.7400 230.4600 54.0200 ;
      RECT 0.0000 52.7400 1.4200 54.0200 ;
      RECT 229.0400 52.3200 229.8350 52.7400 ;
      RECT 0.6250 52.3200 1.4200 52.7400 ;
      RECT 229.0400 51.3800 230.4600 52.3200 ;
      RECT 0.0000 51.3800 1.4200 52.3200 ;
      RECT 229.0400 50.9600 229.8350 51.3800 ;
      RECT 0.6250 50.9600 1.4200 51.3800 ;
      RECT 229.0400 49.6800 230.4600 50.9600 ;
      RECT 0.0000 49.6800 1.4200 50.9600 ;
      RECT 229.0400 49.2600 229.8350 49.6800 ;
      RECT 0.6250 49.2600 1.4200 49.6800 ;
      RECT 229.0400 48.3200 230.4600 49.2600 ;
      RECT 0.0000 48.3200 1.4200 49.2600 ;
      RECT 229.0400 47.9000 229.8350 48.3200 ;
      RECT 0.6250 47.9000 1.4200 48.3200 ;
      RECT 229.0400 46.9600 230.4600 47.9000 ;
      RECT 0.0000 46.9600 1.4200 47.9000 ;
      RECT 229.0400 46.5400 229.8350 46.9600 ;
      RECT 0.6250 46.5400 1.4200 46.9600 ;
      RECT 229.0400 45.2600 230.4600 46.5400 ;
      RECT 0.0000 45.2600 1.4200 46.5400 ;
      RECT 229.0400 44.8400 229.8350 45.2600 ;
      RECT 0.6250 44.8400 1.4200 45.2600 ;
      RECT 229.0400 43.9000 230.4600 44.8400 ;
      RECT 0.0000 43.9000 1.4200 44.8400 ;
      RECT 229.0400 43.4800 229.8350 43.9000 ;
      RECT 0.6250 43.4800 1.4200 43.9000 ;
      RECT 229.0400 42.2000 230.4600 43.4800 ;
      RECT 0.0000 42.2000 1.4200 43.4800 ;
      RECT 229.0400 41.7800 229.8350 42.2000 ;
      RECT 0.6250 41.7800 1.4200 42.2000 ;
      RECT 229.0400 40.8400 230.4600 41.7800 ;
      RECT 0.0000 40.8400 1.4200 41.7800 ;
      RECT 229.0400 40.4200 229.8350 40.8400 ;
      RECT 0.6250 40.4200 1.4200 40.8400 ;
      RECT 229.0400 39.1400 230.4600 40.4200 ;
      RECT 0.0000 39.1400 1.4200 40.4200 ;
      RECT 229.0400 38.7200 229.8350 39.1400 ;
      RECT 0.6250 38.7200 1.4200 39.1400 ;
      RECT 229.0400 37.7800 230.4600 38.7200 ;
      RECT 0.0000 37.7800 1.4200 38.7200 ;
      RECT 229.0400 37.3600 229.8350 37.7800 ;
      RECT 0.6250 37.3600 1.4200 37.7800 ;
      RECT 229.0400 36.4200 230.4600 37.3600 ;
      RECT 0.0000 36.4200 1.4200 37.3600 ;
      RECT 229.0400 36.0000 229.8350 36.4200 ;
      RECT 0.6250 36.0000 1.4200 36.4200 ;
      RECT 229.0400 34.7200 230.4600 36.0000 ;
      RECT 0.0000 34.7200 1.4200 36.0000 ;
      RECT 229.0400 34.3000 229.8350 34.7200 ;
      RECT 0.6250 34.3000 1.4200 34.7200 ;
      RECT 229.0400 33.3600 230.4600 34.3000 ;
      RECT 0.0000 33.3600 1.4200 34.3000 ;
      RECT 229.0400 32.9400 229.8350 33.3600 ;
      RECT 0.6250 32.9400 1.4200 33.3600 ;
      RECT 229.0400 31.6600 230.4600 32.9400 ;
      RECT 0.0000 31.6600 1.4200 32.9400 ;
      RECT 229.0400 31.2400 229.8350 31.6600 ;
      RECT 0.6250 31.2400 1.4200 31.6600 ;
      RECT 229.0400 30.3000 230.4600 31.2400 ;
      RECT 0.0000 30.3000 1.4200 31.2400 ;
      RECT 229.0400 29.8800 229.8350 30.3000 ;
      RECT 0.6250 29.8800 1.4200 30.3000 ;
      RECT 229.0400 28.6000 230.4600 29.8800 ;
      RECT 0.0000 28.6000 1.4200 29.8800 ;
      RECT 229.0400 28.1800 229.8350 28.6000 ;
      RECT 0.6250 28.1800 1.4200 28.6000 ;
      RECT 229.0400 27.2400 230.4600 28.1800 ;
      RECT 0.0000 27.2400 1.4200 28.1800 ;
      RECT 229.0400 26.8200 229.8350 27.2400 ;
      RECT 0.6250 26.8200 1.4200 27.2400 ;
      RECT 229.0400 25.8800 230.4600 26.8200 ;
      RECT 0.0000 25.8800 1.4200 26.8200 ;
      RECT 229.0400 25.4600 229.8350 25.8800 ;
      RECT 0.6250 25.4600 1.4200 25.8800 ;
      RECT 229.0400 24.1800 230.4600 25.4600 ;
      RECT 0.0000 24.1800 1.4200 25.4600 ;
      RECT 229.0400 23.7600 229.8350 24.1800 ;
      RECT 0.6250 23.7600 1.4200 24.1800 ;
      RECT 229.0400 22.8200 230.4600 23.7600 ;
      RECT 0.0000 22.8200 1.4200 23.7600 ;
      RECT 229.0400 22.4000 229.8350 22.8200 ;
      RECT 0.6250 22.4000 1.4200 22.8200 ;
      RECT 229.0400 21.1200 230.4600 22.4000 ;
      RECT 0.0000 21.1200 1.4200 22.4000 ;
      RECT 229.0400 20.7000 229.8350 21.1200 ;
      RECT 0.6250 20.7000 1.4200 21.1200 ;
      RECT 229.0400 19.7600 230.4600 20.7000 ;
      RECT 0.0000 19.7600 1.4200 20.7000 ;
      RECT 229.0400 19.3400 229.8350 19.7600 ;
      RECT 0.6250 19.3400 1.4200 19.7600 ;
      RECT 229.0400 18.0600 230.4600 19.3400 ;
      RECT 0.0000 18.0600 1.4200 19.3400 ;
      RECT 229.0400 17.6400 229.8350 18.0600 ;
      RECT 0.6250 17.6400 1.4200 18.0600 ;
      RECT 229.0400 16.7000 230.4600 17.6400 ;
      RECT 0.0000 16.7000 1.4200 17.6400 ;
      RECT 229.0400 16.2800 229.8350 16.7000 ;
      RECT 0.6250 16.2800 1.4200 16.7000 ;
      RECT 229.0400 15.3400 230.4600 16.2800 ;
      RECT 0.0000 15.3400 1.4200 16.2800 ;
      RECT 229.0400 14.9200 229.8350 15.3400 ;
      RECT 0.6250 14.9200 1.4200 15.3400 ;
      RECT 225.0400 5.2900 225.7600 224.2100 ;
      RECT 195.0600 5.2900 221.7600 224.2100 ;
      RECT 191.8600 5.2900 193.1800 224.2100 ;
      RECT 165.0600 5.2900 189.9800 224.2100 ;
      RECT 161.8600 5.2900 163.1800 224.2100 ;
      RECT 135.0600 5.2900 159.9800 224.2100 ;
      RECT 131.8600 5.2900 133.1800 224.2100 ;
      RECT 105.0600 5.2900 129.9800 224.2100 ;
      RECT 101.8600 5.2900 103.1800 224.2100 ;
      RECT 75.0600 5.2900 99.9800 224.2100 ;
      RECT 71.8600 5.2900 73.1800 224.2100 ;
      RECT 45.0600 5.2900 69.9800 224.2100 ;
      RECT 41.8600 5.2900 43.1800 224.2100 ;
      RECT 15.0600 5.2900 39.9800 224.2100 ;
      RECT 8.7000 5.2900 13.1800 224.2100 ;
      RECT 4.7000 5.2900 5.4200 224.2100 ;
      RECT 229.0400 1.2900 230.4600 14.9200 ;
      RECT 195.0600 1.2900 225.7600 5.2900 ;
      RECT 165.0600 1.2900 193.1800 5.2900 ;
      RECT 135.0600 1.2900 163.1800 5.2900 ;
      RECT 105.0600 1.2900 133.1800 5.2900 ;
      RECT 75.0600 1.2900 103.1800 5.2900 ;
      RECT 45.0600 1.2900 73.1800 5.2900 ;
      RECT 15.0600 1.2900 43.1800 5.2900 ;
      RECT 4.7000 1.2900 13.1800 5.2900 ;
      RECT 0.0000 1.2900 1.4200 14.9200 ;
      RECT 0.0000 0.6250 230.4600 1.2900 ;
      RECT 214.3400 0.0000 230.4600 0.6250 ;
      RECT 209.7400 0.0000 213.9200 0.6250 ;
      RECT 204.6800 0.0000 209.3200 0.6250 ;
      RECT 199.6200 0.0000 204.2600 0.6250 ;
      RECT 194.1000 0.0000 199.2000 0.6250 ;
      RECT 189.9600 0.0000 193.6800 0.6250 ;
      RECT 184.9000 0.0000 189.5400 0.6250 ;
      RECT 179.8400 0.0000 184.4800 0.6250 ;
      RECT 174.7800 0.0000 179.4200 0.6250 ;
      RECT 169.7200 0.0000 174.3600 0.6250 ;
      RECT 165.1200 0.0000 169.3000 0.6250 ;
      RECT 160.0600 0.0000 164.7000 0.6250 ;
      RECT 155.0000 0.0000 159.6400 0.6250 ;
      RECT 149.9400 0.0000 154.5800 0.6250 ;
      RECT 144.4200 0.0000 149.5200 0.6250 ;
      RECT 140.2800 0.0000 144.0000 0.6250 ;
      RECT 135.2200 0.0000 139.8600 0.6250 ;
      RECT 129.7000 0.0000 134.8000 0.6250 ;
      RECT 125.1000 0.0000 129.2800 0.6250 ;
      RECT 120.5000 0.0000 124.6800 0.6250 ;
      RECT 0.0000 0.0000 120.0800 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 228.3700 230.4600 229.8400 ;
      RECT 229.2000 224.7700 230.4600 228.3700 ;
      RECT 0.0000 224.7700 1.2600 228.3700 ;
      RECT 0.0000 224.3700 230.4600 224.7700 ;
      RECT 225.2000 220.7700 230.4600 224.3700 ;
      RECT 0.0000 220.7700 5.2600 224.3700 ;
      RECT 0.0000 8.7300 230.4600 220.7700 ;
      RECT 225.2000 5.1300 230.4600 8.7300 ;
      RECT 0.0000 5.1300 5.2600 8.7300 ;
      RECT 0.0000 4.7300 230.4600 5.1300 ;
      RECT 229.2000 1.1300 230.4600 4.7300 ;
      RECT 0.0000 1.1300 1.2600 4.7300 ;
      RECT 0.0000 0.0000 230.4600 1.1300 ;
  END
END RegFile

END LIBRARY
