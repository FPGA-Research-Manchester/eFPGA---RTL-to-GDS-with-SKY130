// Copyright 2021 University of Manchester
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

module RegFile_ConfigMem (FrameData, FrameStrobe, ConfigBits);
	parameter MaxFramesPerCol = 20;
	parameter FrameBitsPerRow = 32;
	parameter NoConfigBits = 366;
	input [FrameBitsPerRow-1:0] FrameData;
	input [MaxFramesPerCol-1:0] FrameStrobe;
	output [NoConfigBits-1:0] ConfigBits;
	wire [32-1:0] frame0;
	wire [32-1:0] frame1;
	wire [32-1:0] frame2;
	wire [32-1:0] frame3;
	wire [16-1:0] frame4;
	wire [12-1:0] frame5;
	wire [16-1:0] frame6;
	wire [16-1:0] frame7;
	wire [16-1:0] frame8;
	wire [16-1:0] frame9;
	wire [16-1:0] frame10;
	wire [16-1:0] frame11;
	wire [16-1:0] frame12;
	wire [16-1:0] frame13;
	wire [16-1:0] frame14;
	wire [16-1:0] frame15;
	wire [16-1:0] frame16;
	wire [16-1:0] frame17;
	wire [16-1:0] frame18;
	wire [2-1:0] frame19;

//instantiate frame latches
	LHQD1 Inst_frame0_bit31(
	.D(FrameData[31]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[209])
	);

	LHQD1 Inst_frame0_bit30(
	.D(FrameData[30]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[208])
	);

	LHQD1 Inst_frame0_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[207])
	);

	LHQD1 Inst_frame0_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[206])
	);

	LHQD1 Inst_frame0_bit27(
	.D(FrameData[27]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[213])
	);

	LHQD1 Inst_frame0_bit26(
	.D(FrameData[26]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[212])
	);

	LHQD1 Inst_frame0_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[211])
	);

	LHQD1 Inst_frame0_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[210])
	);

	LHQD1 Inst_frame0_bit23(
	.D(FrameData[23]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[217])
	);

	LHQD1 Inst_frame0_bit22(
	.D(FrameData[22]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[216])
	);

	LHQD1 Inst_frame0_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[215])
	);

	LHQD1 Inst_frame0_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[214])
	);

	LHQD1 Inst_frame0_bit19(
	.D(FrameData[19]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[221])
	);

	LHQD1 Inst_frame0_bit18(
	.D(FrameData[18]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[220])
	);

	LHQD1 Inst_frame0_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[219])
	);

	LHQD1 Inst_frame0_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[218])
	);

	LHQD1 Inst_frame0_bit15(
	.D(FrameData[15]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[225])
	);

	LHQD1 Inst_frame0_bit14(
	.D(FrameData[14]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[224])
	);

	LHQD1 Inst_frame0_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[223])
	);

	LHQD1 Inst_frame0_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[222])
	);

	LHQD1 Inst_frame0_bit11(
	.D(FrameData[11]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[229])
	);

	LHQD1 Inst_frame0_bit10(
	.D(FrameData[10]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[228])
	);

	LHQD1 Inst_frame0_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[227])
	);

	LHQD1 Inst_frame0_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[226])
	);

	LHQD1 Inst_frame0_bit7(
	.D(FrameData[7]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[233])
	);

	LHQD1 Inst_frame0_bit6(
	.D(FrameData[6]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[232])
	);

	LHQD1 Inst_frame0_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[231])
	);

	LHQD1 Inst_frame0_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[230])
	);

	LHQD1 Inst_frame0_bit3(
	.D(FrameData[3]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[237])
	);

	LHQD1 Inst_frame0_bit2(
	.D(FrameData[2]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[236])
	);

	LHQD1 Inst_frame0_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[235])
	);

	LHQD1 Inst_frame0_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[0]),
	.Q(ConfigBits[234])
	);

	LHQD1 Inst_frame1_bit31(
	.D(FrameData[31]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[241])
	);

	LHQD1 Inst_frame1_bit30(
	.D(FrameData[30]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[240])
	);

	LHQD1 Inst_frame1_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[239])
	);

	LHQD1 Inst_frame1_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[238])
	);

	LHQD1 Inst_frame1_bit27(
	.D(FrameData[27]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[245])
	);

	LHQD1 Inst_frame1_bit26(
	.D(FrameData[26]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[244])
	);

	LHQD1 Inst_frame1_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[243])
	);

	LHQD1 Inst_frame1_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[242])
	);

	LHQD1 Inst_frame1_bit23(
	.D(FrameData[23]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[249])
	);

	LHQD1 Inst_frame1_bit22(
	.D(FrameData[22]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[248])
	);

	LHQD1 Inst_frame1_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[247])
	);

	LHQD1 Inst_frame1_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[246])
	);

	LHQD1 Inst_frame1_bit19(
	.D(FrameData[19]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[253])
	);

	LHQD1 Inst_frame1_bit18(
	.D(FrameData[18]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[252])
	);

	LHQD1 Inst_frame1_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[251])
	);

	LHQD1 Inst_frame1_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[250])
	);

	LHQD1 Inst_frame1_bit15(
	.D(FrameData[15]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[257])
	);

	LHQD1 Inst_frame1_bit14(
	.D(FrameData[14]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[256])
	);

	LHQD1 Inst_frame1_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[255])
	);

	LHQD1 Inst_frame1_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[254])
	);

	LHQD1 Inst_frame1_bit11(
	.D(FrameData[11]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[261])
	);

	LHQD1 Inst_frame1_bit10(
	.D(FrameData[10]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[260])
	);

	LHQD1 Inst_frame1_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[259])
	);

	LHQD1 Inst_frame1_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[258])
	);

	LHQD1 Inst_frame1_bit7(
	.D(FrameData[7]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[265])
	);

	LHQD1 Inst_frame1_bit6(
	.D(FrameData[6]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[264])
	);

	LHQD1 Inst_frame1_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[263])
	);

	LHQD1 Inst_frame1_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[262])
	);

	LHQD1 Inst_frame1_bit3(
	.D(FrameData[3]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[269])
	);

	LHQD1 Inst_frame1_bit2(
	.D(FrameData[2]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[268])
	);

	LHQD1 Inst_frame1_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[267])
	);

	LHQD1 Inst_frame1_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[1]),
	.Q(ConfigBits[266])
	);

	LHQD1 Inst_frame2_bit31(
	.D(FrameData[31]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[273])
	);

	LHQD1 Inst_frame2_bit30(
	.D(FrameData[30]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[272])
	);

	LHQD1 Inst_frame2_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[271])
	);

	LHQD1 Inst_frame2_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[270])
	);

	LHQD1 Inst_frame2_bit27(
	.D(FrameData[27]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[277])
	);

	LHQD1 Inst_frame2_bit26(
	.D(FrameData[26]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[276])
	);

	LHQD1 Inst_frame2_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[275])
	);

	LHQD1 Inst_frame2_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[274])
	);

	LHQD1 Inst_frame2_bit23(
	.D(FrameData[23]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[281])
	);

	LHQD1 Inst_frame2_bit22(
	.D(FrameData[22]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[280])
	);

	LHQD1 Inst_frame2_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[279])
	);

	LHQD1 Inst_frame2_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[278])
	);

	LHQD1 Inst_frame2_bit19(
	.D(FrameData[19]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[285])
	);

	LHQD1 Inst_frame2_bit18(
	.D(FrameData[18]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[284])
	);

	LHQD1 Inst_frame2_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[283])
	);

	LHQD1 Inst_frame2_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[282])
	);

	LHQD1 Inst_frame2_bit15(
	.D(FrameData[15]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[289])
	);

	LHQD1 Inst_frame2_bit14(
	.D(FrameData[14]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[288])
	);

	LHQD1 Inst_frame2_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[287])
	);

	LHQD1 Inst_frame2_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[286])
	);

	LHQD1 Inst_frame2_bit11(
	.D(FrameData[11]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[293])
	);

	LHQD1 Inst_frame2_bit10(
	.D(FrameData[10]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[292])
	);

	LHQD1 Inst_frame2_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[291])
	);

	LHQD1 Inst_frame2_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[290])
	);

	LHQD1 Inst_frame2_bit7(
	.D(FrameData[7]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[297])
	);

	LHQD1 Inst_frame2_bit6(
	.D(FrameData[6]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[296])
	);

	LHQD1 Inst_frame2_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[295])
	);

	LHQD1 Inst_frame2_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[294])
	);

	LHQD1 Inst_frame2_bit3(
	.D(FrameData[3]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[301])
	);

	LHQD1 Inst_frame2_bit2(
	.D(FrameData[2]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[300])
	);

	LHQD1 Inst_frame2_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[299])
	);

	LHQD1 Inst_frame2_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[2]),
	.Q(ConfigBits[298])
	);

	LHQD1 Inst_frame3_bit31(
	.D(FrameData[31]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[305])
	);

	LHQD1 Inst_frame3_bit30(
	.D(FrameData[30]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[304])
	);

	LHQD1 Inst_frame3_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[303])
	);

	LHQD1 Inst_frame3_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[302])
	);

	LHQD1 Inst_frame3_bit27(
	.D(FrameData[27]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[309])
	);

	LHQD1 Inst_frame3_bit26(
	.D(FrameData[26]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[308])
	);

	LHQD1 Inst_frame3_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[307])
	);

	LHQD1 Inst_frame3_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[306])
	);

	LHQD1 Inst_frame3_bit23(
	.D(FrameData[23]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[313])
	);

	LHQD1 Inst_frame3_bit22(
	.D(FrameData[22]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[312])
	);

	LHQD1 Inst_frame3_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[311])
	);

	LHQD1 Inst_frame3_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[310])
	);

	LHQD1 Inst_frame3_bit19(
	.D(FrameData[19]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[317])
	);

	LHQD1 Inst_frame3_bit18(
	.D(FrameData[18]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[316])
	);

	LHQD1 Inst_frame3_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[315])
	);

	LHQD1 Inst_frame3_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[314])
	);

	LHQD1 Inst_frame3_bit15(
	.D(FrameData[15]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[321])
	);

	LHQD1 Inst_frame3_bit14(
	.D(FrameData[14]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[320])
	);

	LHQD1 Inst_frame3_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[319])
	);

	LHQD1 Inst_frame3_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[318])
	);

	LHQD1 Inst_frame3_bit11(
	.D(FrameData[11]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[325])
	);

	LHQD1 Inst_frame3_bit10(
	.D(FrameData[10]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[324])
	);

	LHQD1 Inst_frame3_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[323])
	);

	LHQD1 Inst_frame3_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[322])
	);

	LHQD1 Inst_frame3_bit7(
	.D(FrameData[7]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[329])
	);

	LHQD1 Inst_frame3_bit6(
	.D(FrameData[6]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[328])
	);

	LHQD1 Inst_frame3_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[327])
	);

	LHQD1 Inst_frame3_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[326])
	);

	LHQD1 Inst_frame3_bit3(
	.D(FrameData[3]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[333])
	);

	LHQD1 Inst_frame3_bit2(
	.D(FrameData[2]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[332])
	);

	LHQD1 Inst_frame3_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[331])
	);

	LHQD1 Inst_frame3_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[3]),
	.Q(ConfigBits[330])
	);

	LHQD1 Inst_frame4_bit31(
	.D(FrameData[31]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[29])
	);

	LHQD1 Inst_frame4_bit30(
	.D(FrameData[30]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[28])
	);

	LHQD1 Inst_frame4_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[27])
	);

	LHQD1 Inst_frame4_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[26])
	);

	LHQD1 Inst_frame4_bit27(
	.D(FrameData[27]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[33])
	);

	LHQD1 Inst_frame4_bit26(
	.D(FrameData[26]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[32])
	);

	LHQD1 Inst_frame4_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[31])
	);

	LHQD1 Inst_frame4_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[30])
	);

	LHQD1 Inst_frame4_bit23(
	.D(FrameData[23]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[61])
	);

	LHQD1 Inst_frame4_bit22(
	.D(FrameData[22]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[60])
	);

	LHQD1 Inst_frame4_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[59])
	);

	LHQD1 Inst_frame4_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[58])
	);

	LHQD1 Inst_frame4_bit19(
	.D(FrameData[19]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[65])
	);

	LHQD1 Inst_frame4_bit18(
	.D(FrameData[18]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[64])
	);

	LHQD1 Inst_frame4_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[63])
	);

	LHQD1 Inst_frame4_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[4]),
	.Q(ConfigBits[62])
	);

	LHQD1 Inst_frame5_bit30(
	.D(FrameData[30]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[84])
	);

	LHQD1 Inst_frame5_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[83])
	);

	LHQD1 Inst_frame5_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[82])
	);

	LHQD1 Inst_frame5_bit26(
	.D(FrameData[26]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[87])
	);

	LHQD1 Inst_frame5_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[86])
	);

	LHQD1 Inst_frame5_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[85])
	);

	LHQD1 Inst_frame5_bit22(
	.D(FrameData[22]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[98])
	);

	LHQD1 Inst_frame5_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[97])
	);

	LHQD1 Inst_frame5_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[96])
	);

	LHQD1 Inst_frame5_bit18(
	.D(FrameData[18]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[109])
	);

	LHQD1 Inst_frame5_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[108])
	);

	LHQD1 Inst_frame5_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[5]),
	.Q(ConfigBits[107])
	);

	LHQD1 Inst_frame6_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[3])
	);

	LHQD1 Inst_frame6_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[2])
	);

	LHQD1 Inst_frame6_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[5])
	);

	LHQD1 Inst_frame6_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[4])
	);

	LHQD1 Inst_frame6_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[7])
	);

	LHQD1 Inst_frame6_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[6])
	);

	LHQD1 Inst_frame6_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[9])
	);

	LHQD1 Inst_frame6_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[8])
	);

	LHQD1 Inst_frame6_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[11])
	);

	LHQD1 Inst_frame6_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[10])
	);

	LHQD1 Inst_frame6_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[13])
	);

	LHQD1 Inst_frame6_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[12])
	);

	LHQD1 Inst_frame6_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[15])
	);

	LHQD1 Inst_frame6_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[14])
	);

	LHQD1 Inst_frame6_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[17])
	);

	LHQD1 Inst_frame6_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[6]),
	.Q(ConfigBits[16])
	);

	LHQD1 Inst_frame7_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[19])
	);

	LHQD1 Inst_frame7_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[18])
	);

	LHQD1 Inst_frame7_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[21])
	);

	LHQD1 Inst_frame7_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[20])
	);

	LHQD1 Inst_frame7_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[23])
	);

	LHQD1 Inst_frame7_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[22])
	);

	LHQD1 Inst_frame7_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[25])
	);

	LHQD1 Inst_frame7_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[24])
	);

	LHQD1 Inst_frame7_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[35])
	);

	LHQD1 Inst_frame7_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[34])
	);

	LHQD1 Inst_frame7_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[37])
	);

	LHQD1 Inst_frame7_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[36])
	);

	LHQD1 Inst_frame7_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[39])
	);

	LHQD1 Inst_frame7_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[38])
	);

	LHQD1 Inst_frame7_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[41])
	);

	LHQD1 Inst_frame7_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[7]),
	.Q(ConfigBits[40])
	);

	LHQD1 Inst_frame8_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[43])
	);

	LHQD1 Inst_frame8_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[42])
	);

	LHQD1 Inst_frame8_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[45])
	);

	LHQD1 Inst_frame8_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[44])
	);

	LHQD1 Inst_frame8_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[47])
	);

	LHQD1 Inst_frame8_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[46])
	);

	LHQD1 Inst_frame8_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[49])
	);

	LHQD1 Inst_frame8_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[48])
	);

	LHQD1 Inst_frame8_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[51])
	);

	LHQD1 Inst_frame8_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[50])
	);

	LHQD1 Inst_frame8_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[53])
	);

	LHQD1 Inst_frame8_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[52])
	);

	LHQD1 Inst_frame8_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[55])
	);

	LHQD1 Inst_frame8_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[54])
	);

	LHQD1 Inst_frame8_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[57])
	);

	LHQD1 Inst_frame8_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[8]),
	.Q(ConfigBits[56])
	);

	LHQD1 Inst_frame9_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[67])
	);

	LHQD1 Inst_frame9_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[66])
	);

	LHQD1 Inst_frame9_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[69])
	);

	LHQD1 Inst_frame9_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[68])
	);

	LHQD1 Inst_frame9_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[71])
	);

	LHQD1 Inst_frame9_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[70])
	);

	LHQD1 Inst_frame9_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[73])
	);

	LHQD1 Inst_frame9_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[72])
	);

	LHQD1 Inst_frame9_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[75])
	);

	LHQD1 Inst_frame9_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[74])
	);

	LHQD1 Inst_frame9_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[77])
	);

	LHQD1 Inst_frame9_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[76])
	);

	LHQD1 Inst_frame9_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[79])
	);

	LHQD1 Inst_frame9_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[78])
	);

	LHQD1 Inst_frame9_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[81])
	);

	LHQD1 Inst_frame9_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[9]),
	.Q(ConfigBits[80])
	);

	LHQD1 Inst_frame10_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[89])
	);

	LHQD1 Inst_frame10_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[88])
	);

	LHQD1 Inst_frame10_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[91])
	);

	LHQD1 Inst_frame10_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[90])
	);

	LHQD1 Inst_frame10_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[93])
	);

	LHQD1 Inst_frame10_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[92])
	);

	LHQD1 Inst_frame10_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[95])
	);

	LHQD1 Inst_frame10_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[94])
	);

	LHQD1 Inst_frame10_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[100])
	);

	LHQD1 Inst_frame10_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[99])
	);

	LHQD1 Inst_frame10_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[102])
	);

	LHQD1 Inst_frame10_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[101])
	);

	LHQD1 Inst_frame10_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[104])
	);

	LHQD1 Inst_frame10_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[103])
	);

	LHQD1 Inst_frame10_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[106])
	);

	LHQD1 Inst_frame10_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[10]),
	.Q(ConfigBits[105])
	);

	LHQD1 Inst_frame11_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[111])
	);

	LHQD1 Inst_frame11_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[110])
	);

	LHQD1 Inst_frame11_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[113])
	);

	LHQD1 Inst_frame11_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[112])
	);

	LHQD1 Inst_frame11_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[115])
	);

	LHQD1 Inst_frame11_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[114])
	);

	LHQD1 Inst_frame11_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[117])
	);

	LHQD1 Inst_frame11_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[116])
	);

	LHQD1 Inst_frame11_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[119])
	);

	LHQD1 Inst_frame11_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[118])
	);

	LHQD1 Inst_frame11_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[121])
	);

	LHQD1 Inst_frame11_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[120])
	);

	LHQD1 Inst_frame11_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[123])
	);

	LHQD1 Inst_frame11_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[122])
	);

	LHQD1 Inst_frame11_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[125])
	);

	LHQD1 Inst_frame11_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[11]),
	.Q(ConfigBits[124])
	);

	LHQD1 Inst_frame12_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[127])
	);

	LHQD1 Inst_frame12_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[126])
	);

	LHQD1 Inst_frame12_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[129])
	);

	LHQD1 Inst_frame12_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[128])
	);

	LHQD1 Inst_frame12_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[131])
	);

	LHQD1 Inst_frame12_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[130])
	);

	LHQD1 Inst_frame12_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[133])
	);

	LHQD1 Inst_frame12_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[132])
	);

	LHQD1 Inst_frame12_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[135])
	);

	LHQD1 Inst_frame12_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[134])
	);

	LHQD1 Inst_frame12_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[137])
	);

	LHQD1 Inst_frame12_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[136])
	);

	LHQD1 Inst_frame12_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[139])
	);

	LHQD1 Inst_frame12_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[138])
	);

	LHQD1 Inst_frame12_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[141])
	);

	LHQD1 Inst_frame12_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[12]),
	.Q(ConfigBits[140])
	);

	LHQD1 Inst_frame13_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[143])
	);

	LHQD1 Inst_frame13_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[142])
	);

	LHQD1 Inst_frame13_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[145])
	);

	LHQD1 Inst_frame13_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[144])
	);

	LHQD1 Inst_frame13_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[147])
	);

	LHQD1 Inst_frame13_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[146])
	);

	LHQD1 Inst_frame13_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[149])
	);

	LHQD1 Inst_frame13_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[148])
	);

	LHQD1 Inst_frame13_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[151])
	);

	LHQD1 Inst_frame13_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[150])
	);

	LHQD1 Inst_frame13_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[153])
	);

	LHQD1 Inst_frame13_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[152])
	);

	LHQD1 Inst_frame13_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[155])
	);

	LHQD1 Inst_frame13_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[154])
	);

	LHQD1 Inst_frame13_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[157])
	);

	LHQD1 Inst_frame13_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[13]),
	.Q(ConfigBits[156])
	);

	LHQD1 Inst_frame14_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[159])
	);

	LHQD1 Inst_frame14_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[158])
	);

	LHQD1 Inst_frame14_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[161])
	);

	LHQD1 Inst_frame14_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[160])
	);

	LHQD1 Inst_frame14_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[163])
	);

	LHQD1 Inst_frame14_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[162])
	);

	LHQD1 Inst_frame14_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[165])
	);

	LHQD1 Inst_frame14_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[164])
	);

	LHQD1 Inst_frame14_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[167])
	);

	LHQD1 Inst_frame14_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[166])
	);

	LHQD1 Inst_frame14_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[169])
	);

	LHQD1 Inst_frame14_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[168])
	);

	LHQD1 Inst_frame14_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[171])
	);

	LHQD1 Inst_frame14_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[170])
	);

	LHQD1 Inst_frame14_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[173])
	);

	LHQD1 Inst_frame14_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[14]),
	.Q(ConfigBits[172])
	);

	LHQD1 Inst_frame15_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[175])
	);

	LHQD1 Inst_frame15_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[174])
	);

	LHQD1 Inst_frame15_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[177])
	);

	LHQD1 Inst_frame15_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[176])
	);

	LHQD1 Inst_frame15_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[179])
	);

	LHQD1 Inst_frame15_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[178])
	);

	LHQD1 Inst_frame15_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[181])
	);

	LHQD1 Inst_frame15_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[180])
	);

	LHQD1 Inst_frame15_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[183])
	);

	LHQD1 Inst_frame15_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[182])
	);

	LHQD1 Inst_frame15_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[185])
	);

	LHQD1 Inst_frame15_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[184])
	);

	LHQD1 Inst_frame15_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[187])
	);

	LHQD1 Inst_frame15_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[186])
	);

	LHQD1 Inst_frame15_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[189])
	);

	LHQD1 Inst_frame15_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[15]),
	.Q(ConfigBits[188])
	);

	LHQD1 Inst_frame16_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[191])
	);

	LHQD1 Inst_frame16_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[190])
	);

	LHQD1 Inst_frame16_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[193])
	);

	LHQD1 Inst_frame16_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[192])
	);

	LHQD1 Inst_frame16_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[195])
	);

	LHQD1 Inst_frame16_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[194])
	);

	LHQD1 Inst_frame16_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[197])
	);

	LHQD1 Inst_frame16_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[196])
	);

	LHQD1 Inst_frame16_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[199])
	);

	LHQD1 Inst_frame16_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[198])
	);

	LHQD1 Inst_frame16_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[201])
	);

	LHQD1 Inst_frame16_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[200])
	);

	LHQD1 Inst_frame16_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[203])
	);

	LHQD1 Inst_frame16_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[202])
	);

	LHQD1 Inst_frame16_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[205])
	);

	LHQD1 Inst_frame16_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[16]),
	.Q(ConfigBits[204])
	);

	LHQD1 Inst_frame17_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[335])
	);

	LHQD1 Inst_frame17_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[334])
	);

	LHQD1 Inst_frame17_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[337])
	);

	LHQD1 Inst_frame17_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[336])
	);

	LHQD1 Inst_frame17_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[339])
	);

	LHQD1 Inst_frame17_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[338])
	);

	LHQD1 Inst_frame17_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[341])
	);

	LHQD1 Inst_frame17_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[340])
	);

	LHQD1 Inst_frame17_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[343])
	);

	LHQD1 Inst_frame17_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[342])
	);

	LHQD1 Inst_frame17_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[345])
	);

	LHQD1 Inst_frame17_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[344])
	);

	LHQD1 Inst_frame17_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[347])
	);

	LHQD1 Inst_frame17_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[346])
	);

	LHQD1 Inst_frame17_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[349])
	);

	LHQD1 Inst_frame17_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[17]),
	.Q(ConfigBits[348])
	);

	LHQD1 Inst_frame18_bit29(
	.D(FrameData[29]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[351])
	);

	LHQD1 Inst_frame18_bit28(
	.D(FrameData[28]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[350])
	);

	LHQD1 Inst_frame18_bit25(
	.D(FrameData[25]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[353])
	);

	LHQD1 Inst_frame18_bit24(
	.D(FrameData[24]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[352])
	);

	LHQD1 Inst_frame18_bit21(
	.D(FrameData[21]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[355])
	);

	LHQD1 Inst_frame18_bit20(
	.D(FrameData[20]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[354])
	);

	LHQD1 Inst_frame18_bit17(
	.D(FrameData[17]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[357])
	);

	LHQD1 Inst_frame18_bit16(
	.D(FrameData[16]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[356])
	);

	LHQD1 Inst_frame18_bit13(
	.D(FrameData[13]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[359])
	);

	LHQD1 Inst_frame18_bit12(
	.D(FrameData[12]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[358])
	);

	LHQD1 Inst_frame18_bit9(
	.D(FrameData[9]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[361])
	);

	LHQD1 Inst_frame18_bit8(
	.D(FrameData[8]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[360])
	);

	LHQD1 Inst_frame18_bit5(
	.D(FrameData[5]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[363])
	);

	LHQD1 Inst_frame18_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[362])
	);

	LHQD1 Inst_frame18_bit1(
	.D(FrameData[1]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[365])
	);

	LHQD1 Inst_frame18_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[18]),
	.Q(ConfigBits[364])
	);

	LHQD1 Inst_frame19_bit4(
	.D(FrameData[4]),
	.E(FrameStrobe[19]),
	.Q(ConfigBits[0])
	);

	LHQD1 Inst_frame19_bit0(
	.D(FrameData[0]),
	.E(FrameStrobe[19]),
	.Q(ConfigBits[1])
	);

endmodule
