##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Wed Apr 21 17:42:26 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO CPU_IO
  CLASS BLOCK ;
  SIZE 29.9000 BY 229.8400 ;
  FOREIGN CPU_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.9924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.844 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.7873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.9731 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 67.4200 0.5950 67.5600 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2655 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.223 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 2.54559 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 9.37239 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 66.0600 0.5950 66.2000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0485 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.101 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 3.05522 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 13.9542 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 64.7000 0.5950 64.8400 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3873 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7915 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.9466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 25.9357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 137.085 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0884848 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 63.0000 0.5950 63.1400 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 79.6600 0.5950 79.8000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0509 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.15 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 3.8369 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 14.936 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 77.9600 0.5950 78.1000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0257 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.061 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 1.67771 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 7.16633 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 76.6000 0.5950 76.7400 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 75.2400 0.5950 75.3800 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 73.5400 0.5950 73.6800 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9061 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3855 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.298 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.27407 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.3805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 72.1800 0.5950 72.3200 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9939 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.398 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4875 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.6316 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 70.4800 0.5950 70.6200 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 69.1200 0.5950 69.2600 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 91.5600 0.5950 91.7000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0509 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.15 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 3.21414 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 14.2034 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 90.2000 0.5950 90.3400 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.55 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.4916 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 88.5000 0.5950 88.6400 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 87.1400 0.5950 87.2800 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 85.7800 0.5950 85.9200 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8605 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 36.0626 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.164 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.0800 0.5950 84.2200 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1185 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 2.34761 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 8.38249 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 82.7200 0.5950 82.8600 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.0000 81.0200 0.5950 81.1600 ;
    END
  END E2END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9915 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.328 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3971 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.5836 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 109.5800 0.5950 109.7200 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1998 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.827 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met1  ;
    ANTENNAMAXAREACAR 10.2388 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 30.9387 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 108.2200 0.5950 108.3600 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6683 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.162 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4261 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.8716 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.265597 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 106.8600 0.5950 107.0000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3346 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.501 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met1  ;
    ANTENNAMAXAREACAR 8.84553 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 23.9725 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 105.1600 0.5950 105.3000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met1  ;
    ANTENNAMAXAREACAR 6.07086 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 20.4758 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 103.8000 0.5950 103.9400 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3315 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.445 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 24.5075 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 97.3651 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 26.313 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 102.1000 0.5950 102.2400 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.043 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.043 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met1  ;
    ANTENNAMAXAREACAR 7.07199 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 26.2642 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 100.7400 0.5950 100.8800 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4281 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.928 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 21.4425 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 96.6905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 22.6347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.462 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 99.0400 0.5950 99.1800 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3285 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.404 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 12.2046 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.1925 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 97.6800 0.5950 97.8200 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2123 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.92 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met1  ;
    ANTENNAMAXAREACAR 5.74763 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.7623 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 96.3200 0.5950 96.4600 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3905 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.48 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.164 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2265 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.302 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 94.6200 0.5950 94.7600 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3369 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.543 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met1  ;
    ANTENNAMAXAREACAR 6.28828 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 21.1655 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 93.2600 0.5950 93.4000 ;
    END
  END E6END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0401 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.8233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.2797 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.616 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 19.4800 0.5950 19.6200 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2609 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 17.7800 0.5950 17.9200 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 16.4200 0.5950 16.5600 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 15.0600 0.5950 15.2000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3701 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.746 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 31.3800 0.5950 31.5200 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8773 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.512 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 30.0200 0.5950 30.1600 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.9778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.352 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 28.3200 0.5950 28.4600 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9445 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 26.9600 0.5950 27.1000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.921 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.4004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.88 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.6000 0.5950 25.7400 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4097 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.464 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 23.9000 0.5950 24.0400 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2133 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.5400 0.5950 22.6800 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6107 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8715 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.304 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 20.8400 0.5950 20.9800 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7685 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.664 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 43.6200 0.5950 43.7600 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.6538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.624 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 41.9200 0.5950 42.0600 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.6766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.216 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 40.5600 0.5950 40.7000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.256 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 38.8600 0.5950 39.0000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.18 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 37.5000 0.5950 37.6400 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5669 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 36.1400 0.5950 36.2800 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6137 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.9132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.448 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 34.4400 0.5950 34.5800 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.4079 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.935 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 32.7400 0.5950 32.8800 ;
    END
  END W2BEGb[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5735 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.61 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 61.6400 0.5950 61.7800 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.6248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 249.136 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 59.9400 0.5950 60.0800 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2931 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.361 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 58.5800 0.5950 58.7200 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7699 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7415 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.88 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 57.2200 0.5950 57.3600 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 55.5200 0.5950 55.6600 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0065 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.1218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.12 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 54.1600 0.5950 54.3000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.2473 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 52.4600 0.5950 52.6000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9865 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.936 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 51.1000 0.5950 51.2400 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.7648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.216 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 49.4000 0.5950 49.5400 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8591 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.452 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 48.0400 0.5950 48.1800 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.1797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.794 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 46.6800 0.5950 46.8200 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.6128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.944 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 44.9800 0.5950 45.1200 ;
    END
  END W6BEG[0]
  PIN OPA_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.239 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 10.4438 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 42.9137 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 105.1600 29.9000 105.3000 ;
    END
  END OPA_I0
  PIN OPA_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6197 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 18.8802 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.3086 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.396701 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 106.5200 29.9000 106.6600 ;
    END
  END OPA_I1
  PIN OPA_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9321 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.485 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 19.6647 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 79.8413 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 24.0684 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.544 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 108.2200 29.9000 108.3600 ;
    END
  END OPA_I2
  PIN OPA_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2625 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.198 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 15.1202 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 67.7939 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.324444 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8867 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.3107 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 109.9200 29.9000 110.0600 ;
    END
  END OPA_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.304 LAYER met4  ;
    ANTENNAMAXAREACAR 3.89646 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 18.8535 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0570313 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 14.8800 0.0000 15.0200 0.4850 ;
    END
  END UserCLK
  PIN OPB_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4947 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.406 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 11.3443 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 28.241 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 98.7000 29.9000 98.8400 ;
    END
  END OPB_I0
  PIN OPB_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2814 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1945 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 32.9639 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 136.139 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.806 LAYER met2  ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 45.3023 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 197.199 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 100.4000 29.9000 100.5400 ;
    END
  END OPB_I1
  PIN OPB_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3966 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.774 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 9.08993 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 34.7355 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 101.7600 29.9000 101.9000 ;
    END
  END OPB_I2
  PIN OPB_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4265 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7049 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.3838 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.293776 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 103.4600 29.9000 103.6000 ;
    END
  END OPB_I3
  PIN RES0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0337 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 92.5800 29.9000 92.7200 ;
    END
  END RES0_O0
  PIN RES0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.7289 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.54 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 93.9400 29.9000 94.0800 ;
    END
  END RES0_O1
  PIN RES0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.6305 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.048 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 95.6400 29.9000 95.7800 ;
    END
  END RES0_O2
  PIN RES0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1268 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5295 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 97.0000 29.9000 97.1400 ;
    END
  END RES0_O3
  PIN RES1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1332 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.558 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3836 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.682 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 86.1200 29.9000 86.2600 ;
    END
  END RES1_O0
  PIN RES1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7901 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.846 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 87.8200 29.9000 87.9600 ;
    END
  END RES1_O1
  PIN RES1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.9525 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.658 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 89.1800 29.9000 89.3200 ;
    END
  END RES1_O2
  PIN RES1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2125 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.995 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 90.8800 29.9000 91.0200 ;
    END
  END RES1_O3
  PIN RES2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.494 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 80.0000 29.9000 80.1400 ;
    END
  END RES2_O0
  PIN RES2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8109 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.464 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 81.3600 29.9000 81.5000 ;
    END
  END RES2_O1
  PIN RES2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.6995 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 83.0600 29.9000 83.2000 ;
    END
  END RES2_O2
  PIN RES2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.368 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 84.4200 29.9000 84.5600 ;
    END
  END RES2_O3
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.0658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.9134 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.387 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 214.8400 0.8000 215.1400 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7336 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.7956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 293.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.1362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.098 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 211.7900 0.8000 212.0900 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.3748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.4085 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 240.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 208.7400 0.8000 209.0400 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.00741 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.5071 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.6900 0.8000 205.9900 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.5651 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.358 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 202.6400 0.8000 202.9400 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.6508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8209 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 199.5900 0.8000 199.8900 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.04 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0176 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 190.329 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 196.5400 0.8000 196.8400 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5846 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 365.281 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 193.4900 0.8000 193.7900 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.0937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.2539 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 190.4400 0.8000 190.7400 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.6858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5566 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.397 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 187.3900 0.8000 187.6900 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.08902 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 23.534 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 184.3400 0.8000 184.6400 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.7523 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.8902 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 181.2900 0.8000 181.5900 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.644 LAYER met3  ;
    ANTENNAMAXAREACAR 21.7956 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.8096 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.670872 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 178.2400 0.8000 178.5400 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 9.14135 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 22.7608 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.25109 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 175.1900 0.8000 175.4900 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 4.2751 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 15.1281 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.101387 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.1400 0.8000 172.4400 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.644 LAYER met3  ;
    ANTENNAMAXAREACAR 5.76139 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 21.6894 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.347601 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 169.0900 0.8000 169.3900 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.5228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.741 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 279.095 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 166.0400 0.8000 166.3400 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 27.1387 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 142.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 162.9900 0.8000 163.2900 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.2342 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.6377 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 159.9400 0.8000 160.2400 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.4118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.5486 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.516 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 156.8900 0.8000 157.1900 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.7108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.803 LAYER met4  ;
    ANTENNAMAXAREACAR 17.589 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 68.1998 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.421579 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 153.8400 0.8000 154.1400 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.803 LAYER met3  ;
    ANTENNAMAXAREACAR 8.59285 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.3821 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.216425 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 150.7900 0.8000 151.0900 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.7206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met4  ;
    ANTENNAMAXAREACAR 50.1396 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 250.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 147.7400 0.8000 148.0400 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.53253 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.4848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.6348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.856 LAYER met4  ;
    ANTENNAGATEAREA 1.0605 LAYER met4  ;
    ANTENNAMAXAREACAR 38.3955 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.492 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 144.6900 0.8000 144.9900 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 3.05172 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 12.3084 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 141.6400 0.8000 141.9400 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.4071 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 82 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 138.5900 0.8000 138.8900 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 32.612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 172.267 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 135.5400 0.8000 135.8400 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.7108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 28.2772 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.879 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 132.4900 0.8000 132.7900 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.803 LAYER met3  ;
    ANTENNAMAXAREACAR 17.1089 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.2561 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.41308 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 129.4400 0.8000 129.7400 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met3  ;
    ANTENNAMAXAREACAR 16.7706 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.1054 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.684259 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 126.3900 0.8000 126.6900 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.803 LAYER met3  ;
    ANTENNAMAXAREACAR 9.57036 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.1115 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.345456 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 123.3400 0.8000 123.6400 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.803 LAYER met3  ;
    ANTENNAMAXAREACAR 7.13129 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.1036 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.345456 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 120.2900 0.8000 120.5900 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1116 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.3056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.904 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 214.8400 29.9000 215.1400 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9069 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.24 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 211.7900 29.9000 212.0900 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 208.7400 29.9000 209.0400 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 205.6900 29.9000 205.9900 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.264 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 202.6400 29.9000 202.9400 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3409 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 199.5900 29.9000 199.8900 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 196.5400 29.9000 196.8400 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.384 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 193.4900 29.9000 193.7900 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.856 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 190.4400 29.9000 190.7400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.76 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 187.3900 29.9000 187.6900 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 184.3400 29.9000 184.6400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 181.2900 29.9000 181.5900 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 178.2400 29.9000 178.5400 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 175.1900 29.9000 175.4900 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 172.1400 29.9000 172.4400 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 169.0900 29.9000 169.3900 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.896 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 166.0400 29.9000 166.3400 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 162.9900 29.9000 163.2900 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 159.9400 29.9000 160.2400 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1706 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.048 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 156.8900 29.9000 157.1900 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.616 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 153.8400 29.9000 154.1400 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 150.7900 29.9000 151.0900 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 147.7400 29.9000 148.0400 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 144.6900 29.9000 144.9900 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 141.6400 29.9000 141.9400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 138.5900 29.9000 138.8900 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 135.5400 29.9000 135.8400 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.5498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.736 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 132.4900 29.9000 132.7900 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.3078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.112 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 129.4400 29.9000 129.7400 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.856 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 126.3900 29.9000 126.6900 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 123.3400 29.9000 123.6400 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 120.2900 29.9000 120.5900 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.3095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.37 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 0.0000 24.6800 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.583 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.8888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 186.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 55.661 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.842 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 22.2400 0.0000 22.3800 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.1495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 29.2572 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.842 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 20.4000 0.0000 20.5400 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.3476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.6007 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 18.5600 0.0000 18.7000 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.4335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9716 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.584 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 16.7200 0.0000 16.8600 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.9576 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 12.5800 0.0000 12.7200 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.179 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.1716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.8749 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.484 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 10.7400 0.0000 10.8800 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.6758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 42.1236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.762 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 8.9000 0.0000 9.0400 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.22 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.3968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7859 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.502 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 7.0600 0.0000 7.2000 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.73306 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.4404 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 5.2200 0.0000 5.3600 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9628 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.696 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met2  ;
    ANTENNAMAXAREACAR 3.79562 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.3414 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0346128 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 0.0000 24.6950 0.3300 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.24 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.126 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 7.17441 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 30.1764 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 0.0000 22.3950 0.3300 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.85859 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.0054 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 19.9250 0.0000 20.0950 0.3300 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.4708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8874 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.752 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 0.0000 18.2550 0.3300 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.694 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.396 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 5.89414 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 25.8586 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 15.7850 0.0000 15.9550 0.3300 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.058 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.011 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 0.0000 13.6550 0.3300 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 12.31 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.432 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.9084 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 11.6450 0.0000 11.8150 0.3300 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.9888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.2593 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 358.498 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 9.3450 0.0000 9.5150 0.3300 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.3309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 24.1884 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.3192 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 25.0123 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.181 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 26.8522 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.171 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.680839 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 7.0450 0.0000 7.2150 0.3300 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.39785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.4752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.022 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6388 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.3089 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.505031 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 0.0000 5.3750 0.3300 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.656 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 229.3550 24.6800 229.8400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.2400 229.3550 22.3800 229.8400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.9400 229.3550 20.0800 229.8400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.1000 229.3550 18.2400 229.8400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.7778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 15.8000 229.3550 15.9400 229.8400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.6978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 13.5000 229.3550 13.6400 229.8400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.294 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 11.6600 229.3550 11.8000 229.8400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.3600 229.3550 9.5000 229.8400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.316 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 7.0600 229.3550 7.2000 229.8400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.9428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 5.2200 229.3550 5.3600 229.8400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.1852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.808 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 229.5100 24.6950 229.8400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.45025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.765 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.242 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 229.5100 22.3950 229.8400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.242 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 19.9250 229.5100 20.0950 229.8400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.462 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 229.5100 18.2550 229.8400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.7850 229.5100 15.9550 229.8400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.2432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.098 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 229.5100 13.6550 229.8400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.8344 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.061 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 11.6450 229.5100 11.8150 229.8400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.06805 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.433 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.268 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 9.3450 229.5100 9.5150 229.8400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.146 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 7.0450 229.5100 7.2150 229.8400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.3756 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.804 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 229.5100 5.3750 229.8400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 24.9100 5.4300 26.4100 224.0700 ;
        RECT 3.4900 5.4300 4.9900 224.0700 ;
      LAYER met3 ;
        RECT 3.4900 5.4300 26.4100 6.9300 ;
        RECT 3.4900 222.5700 26.4100 224.0700 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 27.4100 2.9300 28.9100 226.5700 ;
        RECT 0.9900 2.9300 2.4900 226.5700 ;
      LAYER met3 ;
        RECT 0.9900 2.9300 28.9100 4.4300 ;
        RECT 0.9900 225.0700 28.9100 226.5700 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 24.8650 229.3400 29.9000 229.8400 ;
      RECT 22.5650 229.3400 24.3550 229.8400 ;
      RECT 20.2650 229.3400 22.0550 229.8400 ;
      RECT 18.4250 229.3400 19.7550 229.8400 ;
      RECT 16.1250 229.3400 17.9150 229.8400 ;
      RECT 13.8250 229.3400 15.6150 229.8400 ;
      RECT 11.9850 229.3400 13.3150 229.8400 ;
      RECT 9.6850 229.3400 11.4750 229.8400 ;
      RECT 7.3850 229.3400 9.1750 229.8400 ;
      RECT 5.5450 229.3400 6.8750 229.8400 ;
      RECT 0.0000 229.3400 5.0350 229.8400 ;
      RECT 0.0000 0.5000 29.9000 229.3400 ;
      RECT 24.8650 0.0000 29.9000 0.5000 ;
      RECT 22.5650 0.0000 24.3550 0.5000 ;
      RECT 20.2650 0.0000 22.0550 0.5000 ;
      RECT 18.4250 0.0000 19.7550 0.5000 ;
      RECT 16.1250 0.0000 17.9150 0.5000 ;
      RECT 13.8250 0.0000 15.6150 0.5000 ;
      RECT 11.9850 0.0000 13.3150 0.5000 ;
      RECT 9.6850 0.0000 11.4750 0.5000 ;
      RECT 7.3850 0.0000 9.1750 0.5000 ;
      RECT 5.5450 0.0000 6.8750 0.5000 ;
      RECT 0.0000 0.0000 5.0350 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 110.2000 29.9000 229.8400 ;
      RECT 0.0000 109.8600 29.1650 110.2000 ;
      RECT 0.7350 109.7800 29.1650 109.8600 ;
      RECT 0.7350 109.4400 29.9000 109.7800 ;
      RECT 0.0000 108.5000 29.9000 109.4400 ;
      RECT 0.7350 108.0800 29.1650 108.5000 ;
      RECT 0.0000 107.1400 29.9000 108.0800 ;
      RECT 0.7350 106.8000 29.9000 107.1400 ;
      RECT 0.7350 106.7200 29.1650 106.8000 ;
      RECT 0.0000 106.3800 29.1650 106.7200 ;
      RECT 0.0000 105.4400 29.9000 106.3800 ;
      RECT 0.7350 105.0200 29.1650 105.4400 ;
      RECT 0.0000 104.0800 29.9000 105.0200 ;
      RECT 0.7350 103.7400 29.9000 104.0800 ;
      RECT 0.7350 103.6600 29.1650 103.7400 ;
      RECT 0.0000 103.3200 29.1650 103.6600 ;
      RECT 0.0000 102.3800 29.9000 103.3200 ;
      RECT 0.7350 102.0400 29.9000 102.3800 ;
      RECT 0.7350 101.9600 29.1650 102.0400 ;
      RECT 0.0000 101.6200 29.1650 101.9600 ;
      RECT 0.0000 101.0200 29.9000 101.6200 ;
      RECT 0.7350 100.6800 29.9000 101.0200 ;
      RECT 0.7350 100.6000 29.1650 100.6800 ;
      RECT 0.0000 100.2600 29.1650 100.6000 ;
      RECT 0.0000 99.3200 29.9000 100.2600 ;
      RECT 0.7350 98.9800 29.9000 99.3200 ;
      RECT 0.7350 98.9000 29.1650 98.9800 ;
      RECT 0.0000 98.5600 29.1650 98.9000 ;
      RECT 0.0000 97.9600 29.9000 98.5600 ;
      RECT 0.7350 97.5400 29.9000 97.9600 ;
      RECT 0.0000 97.2800 29.9000 97.5400 ;
      RECT 0.0000 96.8600 29.1650 97.2800 ;
      RECT 0.0000 96.6000 29.9000 96.8600 ;
      RECT 0.7350 96.1800 29.9000 96.6000 ;
      RECT 0.0000 95.9200 29.9000 96.1800 ;
      RECT 0.0000 95.5000 29.1650 95.9200 ;
      RECT 0.0000 94.9000 29.9000 95.5000 ;
      RECT 0.7350 94.4800 29.9000 94.9000 ;
      RECT 0.0000 94.2200 29.9000 94.4800 ;
      RECT 0.0000 93.8000 29.1650 94.2200 ;
      RECT 0.0000 93.5400 29.9000 93.8000 ;
      RECT 0.7350 93.1200 29.9000 93.5400 ;
      RECT 0.0000 92.8600 29.9000 93.1200 ;
      RECT 0.0000 92.4400 29.1650 92.8600 ;
      RECT 0.0000 91.8400 29.9000 92.4400 ;
      RECT 0.7350 91.4200 29.9000 91.8400 ;
      RECT 0.0000 91.1600 29.9000 91.4200 ;
      RECT 0.0000 90.7400 29.1650 91.1600 ;
      RECT 0.0000 90.4800 29.9000 90.7400 ;
      RECT 0.7350 90.0600 29.9000 90.4800 ;
      RECT 0.0000 89.4600 29.9000 90.0600 ;
      RECT 0.0000 89.0400 29.1650 89.4600 ;
      RECT 0.0000 88.7800 29.9000 89.0400 ;
      RECT 0.7350 88.3600 29.9000 88.7800 ;
      RECT 0.0000 88.1000 29.9000 88.3600 ;
      RECT 0.0000 87.6800 29.1650 88.1000 ;
      RECT 0.0000 87.4200 29.9000 87.6800 ;
      RECT 0.7350 87.0000 29.9000 87.4200 ;
      RECT 0.0000 86.4000 29.9000 87.0000 ;
      RECT 0.0000 86.0600 29.1650 86.4000 ;
      RECT 0.7350 85.9800 29.1650 86.0600 ;
      RECT 0.7350 85.6400 29.9000 85.9800 ;
      RECT 0.0000 84.7000 29.9000 85.6400 ;
      RECT 0.0000 84.3600 29.1650 84.7000 ;
      RECT 0.7350 84.2800 29.1650 84.3600 ;
      RECT 0.7350 83.9400 29.9000 84.2800 ;
      RECT 0.0000 83.3400 29.9000 83.9400 ;
      RECT 0.0000 83.0000 29.1650 83.3400 ;
      RECT 0.7350 82.9200 29.1650 83.0000 ;
      RECT 0.7350 82.5800 29.9000 82.9200 ;
      RECT 0.0000 81.6400 29.9000 82.5800 ;
      RECT 0.0000 81.3000 29.1650 81.6400 ;
      RECT 0.7350 81.2200 29.1650 81.3000 ;
      RECT 0.7350 80.8800 29.9000 81.2200 ;
      RECT 0.0000 80.2800 29.9000 80.8800 ;
      RECT 0.0000 79.9400 29.1650 80.2800 ;
      RECT 0.7350 79.8600 29.1650 79.9400 ;
      RECT 0.7350 79.5200 29.9000 79.8600 ;
      RECT 0.0000 78.2400 29.9000 79.5200 ;
      RECT 0.7350 77.8200 29.9000 78.2400 ;
      RECT 0.0000 76.8800 29.9000 77.8200 ;
      RECT 0.7350 76.4600 29.9000 76.8800 ;
      RECT 0.0000 75.5200 29.9000 76.4600 ;
      RECT 0.7350 75.1000 29.9000 75.5200 ;
      RECT 0.0000 73.8200 29.9000 75.1000 ;
      RECT 0.7350 73.4000 29.9000 73.8200 ;
      RECT 0.0000 72.4600 29.9000 73.4000 ;
      RECT 0.7350 72.0400 29.9000 72.4600 ;
      RECT 0.0000 70.7600 29.9000 72.0400 ;
      RECT 0.7350 70.3400 29.9000 70.7600 ;
      RECT 0.0000 69.4000 29.9000 70.3400 ;
      RECT 0.7350 68.9800 29.9000 69.4000 ;
      RECT 0.0000 67.7000 29.9000 68.9800 ;
      RECT 0.7350 67.2800 29.9000 67.7000 ;
      RECT 0.0000 66.3400 29.9000 67.2800 ;
      RECT 0.7350 65.9200 29.9000 66.3400 ;
      RECT 0.0000 64.9800 29.9000 65.9200 ;
      RECT 0.7350 64.5600 29.9000 64.9800 ;
      RECT 0.0000 63.2800 29.9000 64.5600 ;
      RECT 0.7350 62.8600 29.9000 63.2800 ;
      RECT 0.0000 61.9200 29.9000 62.8600 ;
      RECT 0.7350 61.5000 29.9000 61.9200 ;
      RECT 0.0000 60.2200 29.9000 61.5000 ;
      RECT 0.7350 59.8000 29.9000 60.2200 ;
      RECT 0.0000 58.8600 29.9000 59.8000 ;
      RECT 0.7350 58.4400 29.9000 58.8600 ;
      RECT 0.0000 57.5000 29.9000 58.4400 ;
      RECT 0.7350 57.0800 29.9000 57.5000 ;
      RECT 0.0000 55.8000 29.9000 57.0800 ;
      RECT 0.7350 55.3800 29.9000 55.8000 ;
      RECT 0.0000 54.4400 29.9000 55.3800 ;
      RECT 0.7350 54.0200 29.9000 54.4400 ;
      RECT 0.0000 52.7400 29.9000 54.0200 ;
      RECT 0.7350 52.3200 29.9000 52.7400 ;
      RECT 0.0000 51.3800 29.9000 52.3200 ;
      RECT 0.7350 50.9600 29.9000 51.3800 ;
      RECT 0.0000 49.6800 29.9000 50.9600 ;
      RECT 0.7350 49.2600 29.9000 49.6800 ;
      RECT 0.0000 48.3200 29.9000 49.2600 ;
      RECT 0.7350 47.9000 29.9000 48.3200 ;
      RECT 0.0000 46.9600 29.9000 47.9000 ;
      RECT 0.7350 46.5400 29.9000 46.9600 ;
      RECT 0.0000 45.2600 29.9000 46.5400 ;
      RECT 0.7350 44.8400 29.9000 45.2600 ;
      RECT 0.0000 43.9000 29.9000 44.8400 ;
      RECT 0.7350 43.4800 29.9000 43.9000 ;
      RECT 0.0000 42.2000 29.9000 43.4800 ;
      RECT 0.7350 41.7800 29.9000 42.2000 ;
      RECT 0.0000 40.8400 29.9000 41.7800 ;
      RECT 0.7350 40.4200 29.9000 40.8400 ;
      RECT 0.0000 39.1400 29.9000 40.4200 ;
      RECT 0.7350 38.7200 29.9000 39.1400 ;
      RECT 0.0000 37.7800 29.9000 38.7200 ;
      RECT 0.7350 37.3600 29.9000 37.7800 ;
      RECT 0.0000 36.4200 29.9000 37.3600 ;
      RECT 0.7350 36.0000 29.9000 36.4200 ;
      RECT 0.0000 34.7200 29.9000 36.0000 ;
      RECT 0.7350 34.3000 29.9000 34.7200 ;
      RECT 0.0000 33.0200 29.9000 34.3000 ;
      RECT 0.7350 32.6000 29.9000 33.0200 ;
      RECT 0.0000 31.6600 29.9000 32.6000 ;
      RECT 0.7350 31.2400 29.9000 31.6600 ;
      RECT 0.0000 30.3000 29.9000 31.2400 ;
      RECT 0.7350 29.8800 29.9000 30.3000 ;
      RECT 0.0000 28.6000 29.9000 29.8800 ;
      RECT 0.7350 28.1800 29.9000 28.6000 ;
      RECT 0.0000 27.2400 29.9000 28.1800 ;
      RECT 0.7350 26.8200 29.9000 27.2400 ;
      RECT 0.0000 25.8800 29.9000 26.8200 ;
      RECT 0.7350 25.4600 29.9000 25.8800 ;
      RECT 0.0000 24.1800 29.9000 25.4600 ;
      RECT 0.7350 23.7600 29.9000 24.1800 ;
      RECT 0.0000 22.8200 29.9000 23.7600 ;
      RECT 0.7350 22.4000 29.9000 22.8200 ;
      RECT 0.0000 21.1200 29.9000 22.4000 ;
      RECT 0.7350 20.7000 29.9000 21.1200 ;
      RECT 0.0000 19.7600 29.9000 20.7000 ;
      RECT 0.7350 19.3400 29.9000 19.7600 ;
      RECT 0.0000 18.0600 29.9000 19.3400 ;
      RECT 0.7350 17.6400 29.9000 18.0600 ;
      RECT 0.0000 16.7000 29.9000 17.6400 ;
      RECT 0.7350 16.2800 29.9000 16.7000 ;
      RECT 0.0000 15.3400 29.9000 16.2800 ;
      RECT 0.7350 14.9200 29.9000 15.3400 ;
      RECT 0.0000 0.0000 29.9000 14.9200 ;
    LAYER met2 ;
      RECT 24.8200 229.2150 29.9000 229.8400 ;
      RECT 22.5200 229.2150 24.4000 229.8400 ;
      RECT 20.2200 229.2150 22.1000 229.8400 ;
      RECT 18.3800 229.2150 19.8000 229.8400 ;
      RECT 16.0800 229.2150 17.9600 229.8400 ;
      RECT 13.7800 229.2150 15.6600 229.8400 ;
      RECT 11.9400 229.2150 13.3600 229.8400 ;
      RECT 9.6400 229.2150 11.5200 229.8400 ;
      RECT 7.3400 229.2150 9.2200 229.8400 ;
      RECT 5.5000 229.2150 6.9200 229.8400 ;
      RECT 0.0000 229.2150 5.0800 229.8400 ;
      RECT 0.0000 226.7100 29.9000 229.2150 ;
      RECT 2.6300 224.2100 27.2700 226.7100 ;
      RECT 26.5500 5.2900 27.2700 224.2100 ;
      RECT 5.1300 5.2900 24.7700 224.2100 ;
      RECT 2.6300 5.2900 3.3500 224.2100 ;
      RECT 29.0500 2.7900 29.9000 226.7100 ;
      RECT 2.6300 2.7900 27.2700 5.2900 ;
      RECT 0.0000 2.7900 0.8500 226.7100 ;
      RECT 0.0000 0.6250 29.9000 2.7900 ;
      RECT 24.8200 0.0000 29.9000 0.6250 ;
      RECT 22.5200 0.0000 24.4000 0.6250 ;
      RECT 20.6800 0.0000 22.1000 0.6250 ;
      RECT 18.8400 0.0000 20.2600 0.6250 ;
      RECT 17.0000 0.0000 18.4200 0.6250 ;
      RECT 15.1600 0.0000 16.5800 0.6250 ;
      RECT 12.8600 0.0000 14.7400 0.6250 ;
      RECT 11.0200 0.0000 12.4400 0.6250 ;
      RECT 9.1800 0.0000 10.6000 0.6250 ;
      RECT 7.3400 0.0000 8.7600 0.6250 ;
      RECT 5.5000 0.0000 6.9200 0.6250 ;
      RECT 0.0000 0.0000 5.0800 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 226.8700 29.9000 229.8400 ;
      RECT 29.2100 224.7700 29.9000 226.8700 ;
      RECT 0.0000 224.7700 0.6900 226.8700 ;
      RECT 0.0000 224.3700 29.9000 224.7700 ;
      RECT 26.7100 222.2700 29.9000 224.3700 ;
      RECT 0.0000 222.2700 3.1900 224.3700 ;
      RECT 0.0000 215.4400 29.9000 222.2700 ;
      RECT 1.1000 214.5400 28.8000 215.4400 ;
      RECT 0.0000 212.3900 29.9000 214.5400 ;
      RECT 1.1000 211.4900 28.8000 212.3900 ;
      RECT 0.0000 209.3400 29.9000 211.4900 ;
      RECT 1.1000 208.4400 28.8000 209.3400 ;
      RECT 0.0000 206.2900 29.9000 208.4400 ;
      RECT 1.1000 205.3900 28.8000 206.2900 ;
      RECT 0.0000 203.2400 29.9000 205.3900 ;
      RECT 1.1000 202.3400 28.8000 203.2400 ;
      RECT 0.0000 200.1900 29.9000 202.3400 ;
      RECT 1.1000 199.2900 28.8000 200.1900 ;
      RECT 0.0000 197.1400 29.9000 199.2900 ;
      RECT 1.1000 196.2400 28.8000 197.1400 ;
      RECT 0.0000 194.0900 29.9000 196.2400 ;
      RECT 1.1000 193.1900 28.8000 194.0900 ;
      RECT 0.0000 191.0400 29.9000 193.1900 ;
      RECT 1.1000 190.1400 28.8000 191.0400 ;
      RECT 0.0000 187.9900 29.9000 190.1400 ;
      RECT 1.1000 187.0900 28.8000 187.9900 ;
      RECT 0.0000 184.9400 29.9000 187.0900 ;
      RECT 1.1000 184.0400 28.8000 184.9400 ;
      RECT 0.0000 181.8900 29.9000 184.0400 ;
      RECT 1.1000 180.9900 28.8000 181.8900 ;
      RECT 0.0000 178.8400 29.9000 180.9900 ;
      RECT 1.1000 177.9400 28.8000 178.8400 ;
      RECT 0.0000 175.7900 29.9000 177.9400 ;
      RECT 1.1000 174.8900 28.8000 175.7900 ;
      RECT 0.0000 172.7400 29.9000 174.8900 ;
      RECT 1.1000 171.8400 28.8000 172.7400 ;
      RECT 0.0000 169.6900 29.9000 171.8400 ;
      RECT 1.1000 168.7900 28.8000 169.6900 ;
      RECT 0.0000 166.6400 29.9000 168.7900 ;
      RECT 1.1000 165.7400 28.8000 166.6400 ;
      RECT 0.0000 163.5900 29.9000 165.7400 ;
      RECT 1.1000 162.6900 28.8000 163.5900 ;
      RECT 0.0000 160.5400 29.9000 162.6900 ;
      RECT 1.1000 159.6400 28.8000 160.5400 ;
      RECT 0.0000 157.4900 29.9000 159.6400 ;
      RECT 1.1000 156.5900 28.8000 157.4900 ;
      RECT 0.0000 154.4400 29.9000 156.5900 ;
      RECT 1.1000 153.5400 28.8000 154.4400 ;
      RECT 0.0000 151.3900 29.9000 153.5400 ;
      RECT 1.1000 150.4900 28.8000 151.3900 ;
      RECT 0.0000 148.3400 29.9000 150.4900 ;
      RECT 1.1000 147.4400 28.8000 148.3400 ;
      RECT 0.0000 145.2900 29.9000 147.4400 ;
      RECT 1.1000 144.3900 28.8000 145.2900 ;
      RECT 0.0000 142.2400 29.9000 144.3900 ;
      RECT 1.1000 141.3400 28.8000 142.2400 ;
      RECT 0.0000 139.1900 29.9000 141.3400 ;
      RECT 1.1000 138.2900 28.8000 139.1900 ;
      RECT 0.0000 136.1400 29.9000 138.2900 ;
      RECT 1.1000 135.2400 28.8000 136.1400 ;
      RECT 0.0000 133.0900 29.9000 135.2400 ;
      RECT 1.1000 132.1900 28.8000 133.0900 ;
      RECT 0.0000 130.0400 29.9000 132.1900 ;
      RECT 1.1000 129.1400 28.8000 130.0400 ;
      RECT 0.0000 126.9900 29.9000 129.1400 ;
      RECT 1.1000 126.0900 28.8000 126.9900 ;
      RECT 0.0000 123.9400 29.9000 126.0900 ;
      RECT 1.1000 123.0400 28.8000 123.9400 ;
      RECT 0.0000 120.8900 29.9000 123.0400 ;
      RECT 1.1000 119.9900 28.8000 120.8900 ;
      RECT 0.0000 7.2300 29.9000 119.9900 ;
      RECT 26.7100 5.1300 29.9000 7.2300 ;
      RECT 0.0000 5.1300 3.1900 7.2300 ;
      RECT 0.0000 4.7300 29.9000 5.1300 ;
      RECT 29.2100 2.6300 29.9000 4.7300 ;
      RECT 0.0000 2.6300 0.6900 4.7300 ;
      RECT 0.0000 0.0000 29.9000 2.6300 ;
  END
END CPU_IO

END LIBRARY
