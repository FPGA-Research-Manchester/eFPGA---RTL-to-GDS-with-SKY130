##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Thu Apr 22 18:43:40 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO eFPGA_top
  CLASS BLOCK ;
  SIZE 3930.2400 BY 3930.0600 ;
  FOREIGN eFPGA_top 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN I_top[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.107 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3745.2000 0.5950 3745.3400 ;
    END
  END I_top[29]
  PIN I_top[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.0289 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.077 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3733.3000 0.5950 3733.4400 ;
    END
  END I_top[28]
  PIN I_top[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.6553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.209 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3495.3000 0.5950 3495.4400 ;
    END
  END I_top[27]
  PIN I_top[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0725 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.295 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3483.4000 0.5950 3483.5400 ;
    END
  END I_top[26]
  PIN I_top[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.993 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3245.4000 0.5950 3245.5400 ;
    END
  END I_top[25]
  PIN I_top[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0893 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.379 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3233.5000 0.5950 3233.6400 ;
    END
  END I_top[24]
  PIN I_top[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.6217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.041 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2995.5000 0.5950 2995.6400 ;
    END
  END I_top[23]
  PIN I_top[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.1061 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.463 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2983.6000 0.5950 2983.7400 ;
    END
  END I_top[22]
  PIN I_top[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.0289 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.077 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2745.9400 0.5950 2746.0800 ;
    END
  END I_top[21]
  PIN I_top[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0417 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.141 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2733.7000 0.5950 2733.8400 ;
    END
  END I_top[20]
  PIN I_top[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.4085 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.975 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2496.0400 0.5950 2496.1800 ;
    END
  END I_top[19]
  PIN I_top[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.331 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2484.1400 0.5950 2484.2800 ;
    END
  END I_top[18]
  PIN I_top[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.345 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2246.1400 0.5950 2246.2800 ;
    END
  END I_top[17]
  PIN I_top[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.8833 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.349 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2234.2400 0.5950 2234.3800 ;
    END
  END I_top[16]
  PIN I_top[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.107 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1996.2400 0.5950 1996.3800 ;
    END
  END I_top[15]
  PIN I_top[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8869 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.367 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1984.3400 0.5950 1984.4800 ;
    END
  END I_top[14]
  PIN I_top[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0893 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.379 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1746.3400 0.5950 1746.4800 ;
    END
  END I_top[13]
  PIN I_top[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.7273 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.569 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1734.7800 0.5950 1734.9200 ;
    END
  END I_top[12]
  PIN I_top[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.6469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.167 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1496.7800 0.5950 1496.9200 ;
    END
  END I_top[11]
  PIN I_top[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.1849 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.857 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1484.8800 0.5950 1485.0200 ;
    END
  END I_top[10]
  PIN I_top[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.6293 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.079 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1246.8800 0.5950 1247.0200 ;
    END
  END I_top[9]
  PIN I_top[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 12.3241 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.516 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1234.9800 0.5950 1235.1200 ;
    END
  END I_top[8]
  PIN I_top[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.2221 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.043 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 996.9800 0.5950 997.1200 ;
    END
  END I_top[7]
  PIN I_top[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2297 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.044 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 985.0800 0.5950 985.2200 ;
    END
  END I_top[6]
  PIN I_top[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.3273 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.569 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 747.0800 0.5950 747.2200 ;
    END
  END I_top[5]
  PIN I_top[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.1369 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.617 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 735.1800 0.5950 735.3200 ;
    END
  END I_top[4]
  PIN I_top[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.023 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 497.1800 0.5950 497.3200 ;
    END
  END I_top[3]
  PIN I_top[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.8833 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.349 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 485.2800 0.5950 485.4200 ;
    END
  END I_top[2]
  PIN I_top[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.7537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.701 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 247.6200 0.5950 247.7600 ;
    END
  END I_top[1]
  PIN I_top[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8869 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.367 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 235.3800 0.5950 235.5200 ;
    END
  END I_top[0]
  PIN T_top[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.2697 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.281 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3741.1200 0.5950 3741.2600 ;
    END
  END T_top[29]
  PIN T_top[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.107 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3729.2200 0.5950 3729.3600 ;
    END
  END T_top[28]
  PIN T_top[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.9477 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.671 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3491.2200 0.5950 3491.3600 ;
    END
  END T_top[27]
  PIN T_top[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2297 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.044 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3479.3200 0.5950 3479.4600 ;
    END
  END T_top[26]
  PIN T_top[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.331 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3241.3200 0.5950 3241.4600 ;
    END
  END T_top[25]
  PIN T_top[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.9437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.651 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3229.4200 0.5950 3229.5600 ;
    END
  END T_top[24]
  PIN T_top[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.1985 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.925 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2991.4200 0.5950 2991.5600 ;
    END
  END T_top[23]
  PIN T_top[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.0765 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.315 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2979.5200 0.5950 2979.6600 ;
    END
  END T_top[22]
  PIN T_top[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.345 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2741.8600 0.5950 2742.0000 ;
    END
  END T_top[21]
  PIN T_top[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.9437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.651 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2729.9600 0.5950 2730.1000 ;
    END
  END T_top[20]
  PIN T_top[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.3623 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.744 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2491.9600 0.5950 2492.1000 ;
    END
  END T_top[19]
  PIN T_top[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.413 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2480.0600 0.5950 2480.2000 ;
    END
  END T_top[18]
  PIN T_top[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.3777 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.821 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2242.0600 0.5950 2242.2000 ;
    END
  END T_top[17]
  PIN T_top[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.107 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2230.1600 0.5950 2230.3000 ;
    END
  END T_top[16]
  PIN T_top[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8869 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.367 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1992.1600 0.5950 1992.3000 ;
    END
  END T_top[15]
  PIN T_top[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.345 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1980.2600 0.5950 1980.4000 ;
    END
  END T_top[14]
  PIN T_top[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8869 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.367 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1742.2600 0.5950 1742.4000 ;
    END
  END T_top[13]
  PIN T_top[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.345 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1730.3600 0.5950 1730.5000 ;
    END
  END T_top[12]
  PIN T_top[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.6469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.167 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1492.3600 0.5950 1492.5000 ;
    END
  END T_top[11]
  PIN T_top[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.5517 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.691 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1480.8000 0.5950 1480.9400 ;
    END
  END T_top[10]
  PIN T_top[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.4417 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.141 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1242.8000 0.5950 1242.9400 ;
    END
  END T_top[9]
  PIN T_top[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0973 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.419 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1230.9000 0.5950 1231.0400 ;
    END
  END T_top[8]
  PIN T_top[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0417 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.141 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 992.9000 0.5950 993.0400 ;
    END
  END T_top[7]
  PIN T_top[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2657 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.261 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 981.0000 0.5950 981.1400 ;
    END
  END T_top[6]
  PIN T_top[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0893 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.379 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 743.0000 0.5950 743.1400 ;
    END
  END T_top[5]
  PIN T_top[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.345 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 731.1000 0.5950 731.2400 ;
    END
  END T_top[4]
  PIN T_top[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.3301 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.583 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 493.1000 0.5950 493.2400 ;
    END
  END T_top[3]
  PIN T_top[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.107 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 481.2000 0.5950 481.3400 ;
    END
  END T_top[2]
  PIN T_top[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8869 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.367 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 243.2000 0.5950 243.3400 ;
    END
  END T_top[1]
  PIN T_top[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.5265 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.565 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 231.3000 0.5950 231.4400 ;
    END
  END T_top[0]
  PIN O_top[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.878 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 104.181 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.61363 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.1984 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3737.0400 0.5950 3737.1800 ;
    END
  END O_top[29]
  PIN O_top[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9601 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.6555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3725.4800 0.5950 3725.6200 ;
    END
  END O_top[28]
  PIN O_top[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.9648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 104.615 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.62794 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.2699 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3487.1400 0.5950 3487.2800 ;
    END
  END O_top[27]
  PIN O_top[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8565 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.1375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3475.5800 0.5950 3475.7200 ;
    END
  END O_top[26]
  PIN O_top[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.1748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.665 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.66256 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.443 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3237.2400 0.5950 3237.3800 ;
    END
  END O_top[25]
  PIN O_top[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.7809 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.7595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3225.6800 0.5950 3225.8200 ;
    END
  END O_top[24]
  PIN O_top[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.945 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.67179 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.4892 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2987.6800 0.5950 2987.8200 ;
    END
  END O_top[23]
  PIN O_top[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8369 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.0395 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2976.1200 0.5950 2976.2600 ;
    END
  END O_top[22]
  PIN O_top[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.987 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.67317 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.4961 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2737.7800 0.5950 2737.9200 ;
    END
  END O_top[21]
  PIN O_top[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9405 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.5575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2726.2200 0.5950 2726.3600 ;
    END
  END O_top[20]
  PIN O_top[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.074 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.161 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.64594 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.3599 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2487.8800 0.5950 2488.0200 ;
    END
  END O_top[19]
  PIN O_top[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.0441 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.076 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2476.3200 0.5950 2476.4600 ;
    END
  END O_top[18]
  PIN O_top[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.9704 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 104.643 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.62886 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.2746 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2237.9800 0.5950 2238.1200 ;
    END
  END O_top[17]
  PIN O_top[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.1477 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.594 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2226.4200 0.5950 2226.5600 ;
    END
  END O_top[16]
  PIN O_top[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.962 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 104.601 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.62748 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.2676 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1988.0800 0.5950 1988.2200 ;
    END
  END O_top[15]
  PIN O_top[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9489 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.5995 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1976.5200 0.5950 1976.6600 ;
    END
  END O_top[14]
  PIN O_top[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.0488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.035 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.64179 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.3392 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1738.1800 0.5950 1738.3200 ;
    END
  END O_top[13]
  PIN O_top[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.4001 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 101.818 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1726.6200 0.5950 1726.7600 ;
    END
  END O_top[12]
  PIN O_top[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.9648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met3  ;
    ANTENNAMAXAREACAR 9.02899 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 38.3542 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.239668 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1488.6200 0.5950 1488.7600 ;
    END
  END O_top[11]
  PIN O_top[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2333 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.2708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7241 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.6999 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.414531 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1477.0600 0.5950 1477.2000 ;
    END
  END O_top[10]
  PIN O_top[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.3372 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 106.477 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.68933 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.5769 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1238.7200 0.5950 1238.8600 ;
    END
  END O_top[9]
  PIN O_top[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8481 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.0955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1227.1600 0.5950 1227.3000 ;
    END
  END O_top[8]
  PIN O_top[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 106.043 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.67502 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.5053 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 988.8200 0.5950 988.9600 ;
    END
  END O_top[7]
  PIN O_top[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9517 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.6135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 977.2600 0.5950 977.4000 ;
    END
  END O_top[6]
  PIN O_top[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.354 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 106.561 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.6921 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.5907 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 738.9200 0.5950 739.0600 ;
    END
  END O_top[5]
  PIN O_top[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.0553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.132 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 727.3600 0.5950 727.5000 ;
    END
  END O_top[4]
  PIN O_top[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.9592 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 104.587 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.62701 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.2653 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 489.0200 0.5950 489.1600 ;
    END
  END O_top[3]
  PIN O_top[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.0413 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.062 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 477.4600 0.5950 477.6000 ;
    END
  END O_top[2]
  PIN O_top[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.1412 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 105.497 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 5.65702 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 19.4153 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 239.1200 0.5950 239.2600 ;
    END
  END O_top[1]
  PIN O_top[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9377 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.5435 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 1.43396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.09693 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 227.5600 0.5950 227.7000 ;
    END
  END O_top[0]
  PIN OPA[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.7496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.539 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.0489 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 265.939 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3740.1000 3930.2400 3740.2400 ;
    END
  END OPA[59]
  PIN OPA[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5245 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.4775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3741.4600 3930.2400 3741.6000 ;
    END
  END OPA[58]
  PIN OPA[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.8045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0966 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3743.1600 3930.2400 3743.3000 ;
    END
  END OPA[57]
  PIN OPA[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2609 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.302 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3744.8600 3930.2400 3745.0000 ;
    END
  END OPA[56]
  PIN OPA[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.758 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.581 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.0714 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 266.052 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3490.2000 3930.2400 3490.3400 ;
    END
  END OPA[55]
  PIN OPA[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5245 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.4775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.6343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.8825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3491.5600 3930.2400 3491.7000 ;
    END
  END OPA[54]
  PIN OPA[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.918 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 26.5212 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.413 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.76508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3493.2600 3930.2400 3493.4000 ;
    END
  END OPA[53]
  PIN OPA[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.302 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3494.9600 3930.2400 3495.1000 ;
    END
  END OPA[52]
  PIN OPA[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9092 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.337 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.4762 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 268.076 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3240.6400 3930.2400 3240.7800 ;
    END
  END OPA[51]
  PIN OPA[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4845 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.2775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3242.0000 3930.2400 3242.1400 ;
    END
  END OPA[50]
  PIN OPA[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5119 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.4145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 28.7232 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.423 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.76508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3243.7000 3930.2400 3243.8400 ;
    END
  END OPA[49]
  PIN OPA[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.302 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3245.4000 3930.2400 3245.5400 ;
    END
  END OPA[48]
  PIN OPA[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.043 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.3188 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 267.289 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2990.7400 3930.2400 2990.8800 ;
    END
  END OPA[47]
  PIN OPA[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1901 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.8425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2992.1000 3930.2400 2992.2400 ;
    END
  END OPA[46]
  PIN OPA[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3981 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 27.676 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.656 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2993.8000 3930.2400 2993.9400 ;
    END
  END OPA[45]
  PIN OPA[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.9525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 22.5317 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 107.261 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2995.5000 3930.2400 2995.6400 ;
    END
  END OPA[44]
  PIN OPA[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.842 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.001 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.2963 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 267.176 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2740.8400 3930.2400 2740.9800 ;
    END
  END OPA[43]
  PIN OPA[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2769 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.2765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2742.2000 3930.2400 2742.3400 ;
    END
  END OPA[42]
  PIN OPA[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.2665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0966 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2743.9000 3930.2400 2744.0400 ;
    END
  END OPA[41]
  PIN OPA[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4933 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.3585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.4859 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.42 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2745.6000 3930.2400 2745.7400 ;
    END
  END OPA[40]
  PIN OPA[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.435 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.5287 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 268.338 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2490.9400 3930.2400 2491.0800 ;
    END
  END OPA[39]
  PIN OPA[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.6493 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 93.1385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2492.3000 3930.2400 2492.4400 ;
    END
  END OPA[38]
  PIN OPA[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3313 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.5115 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.9498 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.732 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2494.0000 3930.2400 2494.1400 ;
    END
  END OPA[37]
  PIN OPA[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5885 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.8345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0808 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.9247 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.506262 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2495.7000 3930.2400 2495.8400 ;
    END
  END OPA[36]
  PIN OPA[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.73 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.441 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.9964 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 265.677 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2241.0400 3930.2400 2241.1800 ;
    END
  END OPA[35]
  PIN OPA[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5199 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.4175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2242.4000 3930.2400 2242.5400 ;
    END
  END OPA[34]
  PIN OPA[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3621 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.6655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.733 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.553 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2244.1000 3930.2400 2244.2400 ;
    END
  END OPA[33]
  PIN OPA[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4933 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.3585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.5346 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.664 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2245.8000 3930.2400 2245.9400 ;
    END
  END OPA[32]
  PIN OPA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.6656 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.119 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.824 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 264.815 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1991.1400 3930.2400 1991.2800 ;
    END
  END OPA[31]
  PIN OPA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3945 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1992.8400 3930.2400 1992.9800 ;
    END
  END OPA[30]
  PIN OPA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5805 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.7575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0966 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1994.2000 3930.2400 1994.3400 ;
    END
  END OPA[29]
  PIN OPA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1045 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.3775 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.072 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 23.5036 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.039 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.506262 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1995.9000 3930.2400 1996.0400 ;
    END
  END OPA[28]
  PIN OPA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.113 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.3563 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 267.476 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1741.2400 3930.2400 1741.3800 ;
    END
  END OPA[27]
  PIN OPA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.3465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1742.9400 3930.2400 1743.0800 ;
    END
  END OPA[26]
  PIN OPA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4311 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.9735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0966 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1744.3000 3930.2400 1744.4400 ;
    END
  END OPA[25]
  PIN OPA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2497 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.302 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1746.3400 3930.2400 1746.4800 ;
    END
  END OPA[24]
  PIN OPA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.393 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.5062 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 268.226 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1491.6800 3930.2400 1491.8200 ;
    END
  END OPA[23]
  PIN OPA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1873 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.8285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1493.0400 3930.2400 1493.1800 ;
    END
  END OPA[22]
  PIN OPA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4457 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 27.6085 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.319 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1494.7400 3930.2400 1494.8800 ;
    END
  END OPA[21]
  PIN OPA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5885 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.8345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.2546 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 99.4642 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1496.4400 3930.2400 1496.5800 ;
    END
  END OPA[20]
  PIN OPA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.435 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.5287 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 268.338 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1241.7800 3930.2400 1241.9200 ;
    END
  END OPA[19]
  PIN OPA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2685 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.2345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1243.1400 3930.2400 1243.2800 ;
    END
  END OPA[18]
  PIN OPA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3337 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 27.7271 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.324 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1244.8400 3930.2400 1244.9800 ;
    END
  END OPA[17]
  PIN OPA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4765 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.2745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met4  ;
    ANTENNAMAXAREACAR 22.2631 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.194 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.720452 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1246.5400 3930.2400 1246.6800 ;
    END
  END OPA[16]
  PIN OPA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.1276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 100.429 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.0609 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 270.999 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 991.8800 3930.2400 992.0200 ;
    END
  END OPA[15]
  PIN OPA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2769 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.2765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 993.2400 3930.2400 993.3800 ;
    END
  END OPA[14]
  PIN OPA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2637 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.2105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0966 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 994.9400 3930.2400 995.0800 ;
    END
  END OPA[13]
  PIN OPA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4933 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.3585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.376 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 996.6400 3930.2400 996.7800 ;
    END
  END OPA[12]
  PIN OPA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.8224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.903 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 55.2438 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 266.914 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 741.9800 3930.2400 742.1200 ;
    END
  END OPA[11]
  PIN OPA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2853 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.3185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 743.3400 3930.2400 743.4800 ;
    END
  END OPA[10]
  PIN OPA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2077 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.0966 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 745.3800 3930.2400 745.5200 ;
    END
  END OPA[9]
  PIN OPA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4457 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.5271 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.626 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 746.7400 3930.2400 746.8800 ;
    END
  END OPA[8]
  PIN OPA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.7188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.385 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.9664 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 265.527 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 492.0800 3930.2400 492.2200 ;
    END
  END OPA[7]
  PIN OPA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4393 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.0885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 493.4400 3930.2400 493.5800 ;
    END
  END OPA[6]
  PIN OPA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4601 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.786 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 28.2336 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.681 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.76508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 495.1400 3930.2400 495.2800 ;
    END
  END OPA[5]
  PIN OPA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6053 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.9185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.051 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0883 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.9622 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.506262 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 496.8400 3930.2400 496.9800 ;
    END
  END OPA[4]
  PIN OPA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.6628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 98.105 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.8165 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 264.777 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 242.5200 3930.2400 242.6600 ;
    END
  END OPA[3]
  PIN OPA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3833 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.8085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 3.64337 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.6908 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 243.8800 3930.2400 244.0200 ;
    END
  END OPA[2]
  PIN OPA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5861 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.7855 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.786 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 28.5527 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.57 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.76508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 245.5800 3930.2400 245.7200 ;
    END
  END OPA[1]
  PIN OPA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2525 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 21.9552 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 103.302 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.613357 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 247.2800 3930.2400 247.4200 ;
    END
  END OPA[0]
  PIN OPB[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.3095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9711 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.0322 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.137617 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3733.6400 3930.2400 3733.7800 ;
    END
  END OPB[59]
  PIN OPB[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4289 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.0365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.792 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3735.3400 3930.2400 3735.4800 ;
    END
  END OPB[58]
  PIN OPB[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.6315 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1282 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.5842 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3736.7000 3930.2400 3736.8400 ;
    END
  END OPB[57]
  PIN OPB[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.11 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.196 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 28.1598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.026 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.293776 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3738.4000 3930.2400 3738.5400 ;
    END
  END OPB[56]
  PIN OPB[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.9449 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.5795 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.1218 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.7858 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.137617 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3483.7400 3930.2400 3483.8800 ;
    END
  END OPB[55]
  PIN OPB[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5717 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.7505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.95 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3485.4400 3930.2400 3485.5800 ;
    END
  END OPB[54]
  PIN OPB[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.065 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.116 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 53.7175 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 257.873 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3486.8000 3930.2400 3486.9400 ;
    END
  END OPB[53]
  PIN OPB[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.979 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 28.0436 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.445 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.293776 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3488.5000 3930.2400 3488.6400 ;
    END
  END OPB[52]
  PIN OPB[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7381 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.5825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.0248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 66.0372 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 319.66 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.244712 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3234.1800 3930.2400 3234.3200 ;
    END
  END OPB[51]
  PIN OPB[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6277 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.0305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.95 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3235.8800 3930.2400 3236.0200 ;
    END
  END OPB[50]
  PIN OPB[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1658 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.62 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 53.9874 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 259.223 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3237.2400 3930.2400 3237.3800 ;
    END
  END OPB[49]
  PIN OPB[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4331 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.9835 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3238.9400 3930.2400 3239.0800 ;
    END
  END OPB[48]
  PIN OPB[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7733 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7215 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.7868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 83.476 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 412.487 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.244712 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2984.2800 3930.2400 2984.4200 ;
    END
  END OPB[47]
  PIN OPB[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5073 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.4285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.9594 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.171 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2985.9800 3930.2400 2986.1200 ;
    END
  END OPB[46]
  PIN OPB[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1294 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.438 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 53.8899 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 258.736 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2987.3400 3930.2400 2987.4800 ;
    END
  END OPB[45]
  PIN OPB[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9969 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.8765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2989.0400 3930.2400 2989.1800 ;
    END
  END OPB[44]
  PIN OPB[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2359 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.112 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.1668 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 252.353 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2734.3800 3930.2400 2734.5200 ;
    END
  END OPB[43]
  PIN OPB[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.7905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.95 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2736.0800 3930.2400 2736.2200 ;
    END
  END OPB[42]
  PIN OPB[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2442 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.012 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.1973 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 260.272 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2737.4400 3930.2400 2737.5800 ;
    END
  END OPB[41]
  PIN OPB[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1789 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.7865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2739.1400 3930.2400 2739.2800 ;
    END
  END OPB[40]
  PIN OPB[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3333 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.525 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.4276 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 253.459 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2484.4800 3930.2400 2484.6200 ;
    END
  END OPB[39]
  PIN OPB[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4457 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 48.8199 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 215.862 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2486.1800 3930.2400 2486.3200 ;
    END
  END OPB[38]
  PIN OPB[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2358 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.97 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.1748 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 260.16 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2487.5400 3930.2400 2487.6800 ;
    END
  END OPB[37]
  PIN OPB[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.5513 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.6485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2489.2400 3930.2400 2489.3800 ;
    END
  END OPB[36]
  PIN OPB[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2367 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.042 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.1689 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 252.166 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2234.5800 3930.2400 2234.7200 ;
    END
  END OPB[35]
  PIN OPB[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4601 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.0254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.773 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 48.3736 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 212.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.76508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2236.2800 3930.2400 2236.4200 ;
    END
  END OPB[34]
  PIN OPB[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.4402 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.992 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.7221 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 262.896 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2237.6400 3930.2400 2237.7800 ;
    END
  END OPB[33]
  PIN OPB[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2567 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.1015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2239.3400 3930.2400 2239.4800 ;
    END
  END OPB[32]
  PIN OPB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 149.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met4  ;
    ANTENNAMAXAREACAR 18.7531 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 69.7216 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.351807 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1984.6800 3930.2400 1984.8200 ;
    END
  END OPB[31]
  PIN OPB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5885 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.8345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.1422 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 217.473 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1986.7200 3930.2400 1986.8600 ;
    END
  END OPB[30]
  PIN OPB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.481 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.4881 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 261.528 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1987.7400 3930.2400 1987.8800 ;
    END
  END OPB[29]
  PIN OPB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2013 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1989.7800 3930.2400 1989.9200 ;
    END
  END OPB[28]
  PIN OPB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2611 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.238 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.2343 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 252.691 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1735.1200 3930.2400 1735.2600 ;
    END
  END OPB[27]
  PIN OPB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5269 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 47.89 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 209.742 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.76508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1736.8200 3930.2400 1736.9600 ;
    END
  END OPB[26]
  PIN OPB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.0678 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.13 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 53.725 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 257.911 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1738.1800 3930.2400 1738.3200 ;
    END
  END OPB[25]
  PIN OPB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0977 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.3805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1739.8800 3930.2400 1740.0200 ;
    END
  END OPB[24]
  PIN OPB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4901 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.309 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.8474 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 255.558 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1485.2200 3930.2400 1485.3600 ;
    END
  END OPB[23]
  PIN OPB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6053 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.9185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 48.4879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 214.078 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1486.9200 3930.2400 1487.0600 ;
    END
  END OPB[22]
  PIN OPB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1322 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.452 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 53.8974 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 258.773 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1488.2800 3930.2400 1488.4200 ;
    END
  END OPB[21]
  PIN OPB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9941 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.8625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1489.9800 3930.2400 1490.1200 ;
    END
  END OPB[20]
  PIN OPB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0265 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.3008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 66.1427 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 320.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.244712 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1235.3200 3930.2400 1235.4600 ;
    END
  END OPB[19]
  PIN OPB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2721 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.2525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.95 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1237.0200 3930.2400 1237.1600 ;
    END
  END OPB[18]
  PIN OPB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8805 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.2575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9499 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.6927 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1238.3800 3930.2400 1238.5200 ;
    END
  END OPB[17]
  PIN OPB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0809 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.2965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1240.0800 3930.2400 1240.2200 ;
    END
  END OPB[16]
  PIN OPB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4257 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.987 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.675 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 254.696 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 985.4200 3930.2400 985.5600 ;
    END
  END OPB[15]
  PIN OPB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2861 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3594 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.358 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 987.1200 3930.2400 987.2600 ;
    END
  END OPB[14]
  PIN OPB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2912 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.173 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.3231 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 260.703 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 988.4800 3930.2400 988.6200 ;
    END
  END OPB[13]
  PIN OPB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2623 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.1295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 990.1800 3930.2400 990.3200 ;
    END
  END OPB[12]
  PIN OPB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3507 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.686 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.4742 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 253.89 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 735.5200 3930.2400 735.6600 ;
    END
  END OPB[11]
  PIN OPB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2669 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.9631 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.19 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 737.2200 3930.2400 737.3600 ;
    END
  END OPB[10]
  PIN OPB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3478 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 96.53 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 54.4747 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 261.659 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 738.5800 3930.2400 738.7200 ;
    END
  END OPB[9]
  PIN OPB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.0921 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 90.3525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 740.2800 3930.2400 740.4200 ;
    END
  END OPB[8]
  PIN OPB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4543 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.204 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met1  ;
    ANTENNAMAXAREACAR 56.7515 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 255.277 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0773762 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 485.6200 3930.2400 485.7600 ;
    END
  END OPB[7]
  PIN OPB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6669 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.2265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3149 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.136 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 487.3200 3930.2400 487.4600 ;
    END
  END OPB[6]
  PIN OPB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6197 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.9535 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.03 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8996 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.441 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 488.6800 3930.2400 488.8200 ;
    END
  END OPB[5]
  PIN OPB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3413 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.5985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 490.3800 3930.2400 490.5200 ;
    END
  END OPB[4]
  PIN OPB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.001 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met4  ;
    ANTENNAMAXAREACAR 18.0966 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 66.4713 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.351807 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 235.7200 3930.2400 235.8600 ;
    END
  END OPB[3]
  PIN OPB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6669 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.2265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.95 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.872175 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 237.7600 3930.2400 237.9000 ;
    END
  END OPB[2]
  PIN OPB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.3095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1507 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.6967 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.289606 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 238.7800 3930.2400 238.9200 ;
    END
  END OPB[1]
  PIN OPB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2853 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.3185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.98 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5813 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5904 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 240.8200 3930.2400 240.9600 ;
    END
  END OPB[0]
  PIN RES0[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.8361 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.113 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3727.5200 3930.2400 3727.6600 ;
    END
  END RES0[59]
  PIN RES0[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0529 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.197 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3728.8800 3930.2400 3729.0200 ;
    END
  END RES0[58]
  PIN RES0[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0361 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.113 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3730.5800 3930.2400 3730.7200 ;
    END
  END RES0[57]
  PIN RES0[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.447 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3731.9400 3930.2400 3732.0800 ;
    END
  END RES0[56]
  PIN RES0[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.7613 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.739 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3477.6200 3930.2400 3477.7600 ;
    END
  END RES0[55]
  PIN RES0[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8625 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.245 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3478.9800 3930.2400 3479.1200 ;
    END
  END RES0[54]
  PIN RES0[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6325 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.095 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3480.6800 3930.2400 3480.8200 ;
    END
  END RES0[53]
  PIN RES0[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.7037 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.451 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3482.0400 3930.2400 3482.1800 ;
    END
  END RES0[52]
  PIN RES0[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3228.0600 3930.2400 3228.2000 ;
    END
  END RES0[51]
  PIN RES0[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3229.0800 3930.2400 3229.2200 ;
    END
  END RES0[50]
  PIN RES0[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2153 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.009 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3231.1200 3930.2400 3231.2600 ;
    END
  END RES0[49]
  PIN RES0[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9835 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.813 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3232.1400 3930.2400 3232.2800 ;
    END
  END RES0[48]
  PIN RES0[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2978.1600 3930.2400 2978.3000 ;
    END
  END RES0[47]
  PIN RES0[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.792 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2979.5200 3930.2400 2979.6600 ;
    END
  END RES0[46]
  PIN RES0[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.447 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2981.2200 3930.2400 2981.3600 ;
    END
  END RES0[45]
  PIN RES0[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.2257 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.061 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2982.5800 3930.2400 2982.7200 ;
    END
  END RES0[44]
  PIN RES0[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0865 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.365 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2728.2600 3930.2400 2728.4000 ;
    END
  END RES0[43]
  PIN RES0[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0529 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.197 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2729.6200 3930.2400 2729.7600 ;
    END
  END RES0[42]
  PIN RES0[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.9241 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2731.3200 3930.2400 2731.4600 ;
    END
  END RES0[41]
  PIN RES0[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.1921 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.893 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2732.6800 3930.2400 2732.8200 ;
    END
  END RES0[40]
  PIN RES0[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.5001 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.433 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2478.3600 3930.2400 2478.5000 ;
    END
  END RES0[39]
  PIN RES0[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2479.7200 3930.2400 2479.8600 ;
    END
  END RES0[38]
  PIN RES0[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.1921 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.893 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2481.4200 3930.2400 2481.5600 ;
    END
  END RES0[37]
  PIN RES0[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.769 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2482.7800 3930.2400 2482.9200 ;
    END
  END RES0[36]
  PIN RES0[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.1657 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.724 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2228.4600 3930.2400 2228.6000 ;
    END
  END RES0[35]
  PIN RES0[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1817 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.841 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2229.8200 3930.2400 2229.9600 ;
    END
  END RES0[34]
  PIN RES0[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.2597 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.231 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2231.5200 3930.2400 2231.6600 ;
    END
  END RES0[33]
  PIN RES0[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2232.8800 3930.2400 2233.0200 ;
    END
  END RES0[32]
  PIN RES0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9173 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.519 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1978.5600 3930.2400 1978.7000 ;
    END
  END RES0[31]
  PIN RES0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6661 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.263 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1979.9200 3930.2400 1980.0600 ;
    END
  END RES0[30]
  PIN RES0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.7753 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.809 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1981.6200 3930.2400 1981.7600 ;
    END
  END RES0[29]
  PIN RES0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.3227 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.509 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1982.9800 3930.2400 1983.1200 ;
    END
  END RES0[28]
  PIN RES0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1729.0000 3930.2400 1729.1400 ;
    END
  END RES0[27]
  PIN RES0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2129 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.96 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1730.3600 3930.2400 1730.5000 ;
    END
  END RES0[26]
  PIN RES0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3105 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.485 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1732.0600 3930.2400 1732.2000 ;
    END
  END RES0[25]
  PIN RES0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.1757 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.774 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1733.4200 3930.2400 1733.5600 ;
    END
  END RES0[24]
  PIN RES0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1479.1000 3930.2400 1479.2400 ;
    END
  END RES0[23]
  PIN RES0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4701 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.283 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1480.4600 3930.2400 1480.6000 ;
    END
  END RES0[22]
  PIN RES0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.1785 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.825 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1482.1600 3930.2400 1482.3000 ;
    END
  END RES0[21]
  PIN RES0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6801 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.333 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1483.5200 3930.2400 1483.6600 ;
    END
  END RES0[20]
  PIN RES0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.331 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1229.2000 3930.2400 1229.3400 ;
    END
  END RES0[19]
  PIN RES0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.1273 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.569 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1230.5600 3930.2400 1230.7000 ;
    END
  END RES0[18]
  PIN RES0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.329 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1232.2600 3930.2400 1232.4000 ;
    END
  END RES0[17]
  PIN RES0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.5281 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.536 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1233.6200 3930.2400 1233.7600 ;
    END
  END RES0[16]
  PIN RES0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.9889 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.84 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 979.3000 3930.2400 979.4400 ;
    END
  END RES0[15]
  PIN RES0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9341 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.603 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 980.6600 3930.2400 980.8000 ;
    END
  END RES0[14]
  PIN RES0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.3405 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.635 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 982.3600 3930.2400 982.5000 ;
    END
  END RES0[13]
  PIN RES0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.4493 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.179 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 983.7200 3930.2400 983.8600 ;
    END
  END RES0[12]
  PIN RES0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 729.4000 3930.2400 729.5400 ;
    END
  END RES0[11]
  PIN RES0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.1245 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.555 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 730.7600 3930.2400 730.9000 ;
    END
  END RES0[10]
  PIN RES0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.3657 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.724 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 732.4600 3930.2400 732.6000 ;
    END
  END RES0[9]
  PIN RES0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.769 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 733.8200 3930.2400 733.9600 ;
    END
  END RES0[8]
  PIN RES0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3717 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.791 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 479.5000 3930.2400 479.6400 ;
    END
  END RES0[7]
  PIN RES0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.2085 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.975 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 481.2000 3930.2400 481.3400 ;
    END
  END RES0[6]
  PIN RES0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.3689 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.74 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 482.5600 3930.2400 482.7000 ;
    END
  END RES0[5]
  PIN RES0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.6121 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.993 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 484.2600 3930.2400 484.4000 ;
    END
  END RES0[4]
  PIN RES0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1005 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.435 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 229.9400 3930.2400 230.0800 ;
    END
  END RES0[3]
  PIN RES0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3745 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.805 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 231.3000 3930.2400 231.4400 ;
    END
  END RES0[2]
  PIN RES0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.5985 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.925 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 233.0000 3930.2400 233.1400 ;
    END
  END RES0[1]
  PIN RES0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.0461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 234.3600 3930.2400 234.5000 ;
    END
  END RES0[0]
  PIN RES1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.447 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3721.0600 3930.2400 3721.2000 ;
    END
  END RES1[59]
  PIN RES1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.7409 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.637 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3722.7600 3930.2400 3722.9000 ;
    END
  END RES1[58]
  PIN RES1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.331 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3724.1200 3930.2400 3724.2600 ;
    END
  END RES1[57]
  PIN RES1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3725.8200 3930.2400 3725.9600 ;
    END
  END RES1[56]
  PIN RES1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3105 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.485 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3471.1600 3930.2400 3471.3000 ;
    END
  END RES1[55]
  PIN RES1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.7273 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.569 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3472.8600 3930.2400 3473.0000 ;
    END
  END RES1[54]
  PIN RES1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0497 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.181 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3474.2200 3930.2400 3474.3600 ;
    END
  END RES1[53]
  PIN RES1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9509 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.687 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3475.9200 3930.2400 3476.0600 ;
    END
  END RES1[52]
  PIN RES1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6325 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.095 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3221.6000 3930.2400 3221.7400 ;
    END
  END RES1[51]
  PIN RES1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7197 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.531 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3222.9600 3930.2400 3223.1000 ;
    END
  END RES1[50]
  PIN RES1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9341 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.603 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3224.6600 3930.2400 3224.8000 ;
    END
  END RES1[49]
  PIN RES1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.331 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3226.0200 3930.2400 3226.1600 ;
    END
  END RES1[48]
  PIN RES1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.1581 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.723 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2971.7000 3930.2400 2971.8400 ;
    END
  END RES1[47]
  PIN RES1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.9545 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.705 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2973.4000 3930.2400 2973.5400 ;
    END
  END RES1[46]
  PIN RES1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.5309 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.587 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2974.7600 3930.2400 2974.9000 ;
    END
  END RES1[45]
  PIN RES1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3413 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.639 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2976.4600 3930.2400 2976.6000 ;
    END
  END RES1[44]
  PIN RES1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9957 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.911 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2721.8000 3930.2400 2721.9400 ;
    END
  END RES1[43]
  PIN RES1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3105 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.485 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2723.5000 3930.2400 2723.6400 ;
    END
  END RES1[42]
  PIN RES1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7197 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.531 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2724.8600 3930.2400 2725.0000 ;
    END
  END RES1[41]
  PIN RES1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.2085 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.975 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2726.5600 3930.2400 2726.7000 ;
    END
  END RES1[40]
  PIN RES1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8149 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.007 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2471.9000 3930.2400 2472.0400 ;
    END
  END RES1[39]
  PIN RES1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6465 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.165 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2473.6000 3930.2400 2473.7400 ;
    END
  END RES1[38]
  PIN RES1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3441 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.653 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2474.9600 3930.2400 2475.1000 ;
    END
  END RES1[37]
  PIN RES1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3105 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.485 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2476.6600 3930.2400 2476.8000 ;
    END
  END RES1[36]
  PIN RES1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4085 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.975 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2222.0000 3930.2400 2222.1400 ;
    END
  END RES1[35]
  PIN RES1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2223.7000 3930.2400 2223.8400 ;
    END
  END RES1[34]
  PIN RES1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.7409 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.637 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2225.0600 3930.2400 2225.2000 ;
    END
  END RES1[33]
  PIN RES1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.4625 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.245 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2226.7600 3930.2400 2226.9000 ;
    END
  END RES1[32]
  PIN RES1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0865 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.365 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1972.1000 3930.2400 1972.2400 ;
    END
  END RES1[31]
  PIN RES1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.4709 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.25 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1973.8000 3930.2400 1973.9400 ;
    END
  END RES1[30]
  PIN RES1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8741 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.266 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1975.1600 3930.2400 1975.3000 ;
    END
  END RES1[29]
  PIN RES1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4393 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.129 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1976.8600 3930.2400 1977.0000 ;
    END
  END RES1[28]
  PIN RES1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1722.5400 3930.2400 1722.6800 ;
    END
  END RES1[27]
  PIN RES1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.9885 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.875 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1724.2400 3930.2400 1724.3800 ;
    END
  END RES1[26]
  PIN RES1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.6937 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.401 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1725.6000 3930.2400 1725.7400 ;
    END
  END RES1[25]
  PIN RES1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0361 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.113 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1727.3000 3930.2400 1727.4400 ;
    END
  END RES1[24]
  PIN RES1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.2729 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.297 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1472.6400 3930.2400 1472.7800 ;
    END
  END RES1[23]
  PIN RES1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0021 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.943 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1474.3400 3930.2400 1474.4800 ;
    END
  END RES1[22]
  PIN RES1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.8089 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.977 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1475.7000 3930.2400 1475.8400 ;
    END
  END RES1[21]
  PIN RES1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7981 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.923 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1477.4000 3930.2400 1477.5400 ;
    END
  END RES1[20]
  PIN RES1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3717 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.791 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1222.7400 3930.2400 1222.8800 ;
    END
  END RES1[19]
  PIN RES1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6325 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.095 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1224.4400 3930.2400 1224.5800 ;
    END
  END RES1[18]
  PIN RES1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0329 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.097 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1225.8000 3930.2400 1225.9400 ;
    END
  END RES1[17]
  PIN RES1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.3205 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.535 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1227.5000 3930.2400 1227.6400 ;
    END
  END RES1[16]
  PIN RES1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.8697 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.281 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 972.8400 3930.2400 972.9800 ;
    END
  END RES1[15]
  PIN RES1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4533 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.199 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 974.5400 3930.2400 974.6800 ;
    END
  END RES1[14]
  PIN RES1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4393 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.129 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 975.9000 3930.2400 976.0400 ;
    END
  END RES1[13]
  PIN RES1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.9041 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.453 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 977.6000 3930.2400 977.7400 ;
    END
  END RES1[12]
  PIN RES1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.447 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 722.9400 3930.2400 723.0800 ;
    END
  END RES1[11]
  PIN RES1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 724.6400 3930.2400 724.7800 ;
    END
  END RES1[10]
  PIN RES1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2153 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.009 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 726.0000 3930.2400 726.1400 ;
    END
  END RES1[9]
  PIN RES1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.0293 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.079 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 727.7000 3930.2400 727.8400 ;
    END
  END RES1[8]
  PIN RES1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0833 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.349 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 473.0400 3930.2400 473.1800 ;
    END
  END RES1[7]
  PIN RES1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.0769 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.317 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 475.0800 3930.2400 475.2200 ;
    END
  END RES1[6]
  PIN RES1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4729 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.297 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 476.1000 3930.2400 476.2400 ;
    END
  END RES1[5]
  PIN RES1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3409 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.637 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 478.1400 3930.2400 478.2800 ;
    END
  END RES1[4]
  PIN RES1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1173 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.519 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 223.4800 3930.2400 223.6200 ;
    END
  END RES1[3]
  PIN RES1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 11.0217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.041 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 225.1800 3930.2400 225.3200 ;
    END
  END RES1[2]
  PIN RES1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.02 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.0325 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 226.5400 3930.2400 226.6800 ;
    END
  END RES1[1]
  PIN RES1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 228.2400 3930.2400 228.3800 ;
    END
  END RES1[0]
  PIN RES2[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.1921 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.893 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3714.9400 3930.2400 3715.0800 ;
    END
  END RES2[59]
  PIN RES2[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3917 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.891 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3716.3000 3930.2400 3716.4400 ;
    END
  END RES2[58]
  PIN RES2[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.8221 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.043 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3718.0000 3930.2400 3718.1400 ;
    END
  END RES2[57]
  PIN RES2[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5681 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.773 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3719.3600 3930.2400 3719.5000 ;
    END
  END RES2[56]
  PIN RES2[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8561 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.213 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3465.3800 3930.2400 3465.5200 ;
    END
  END RES2[55]
  PIN RES2[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.8337 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.064 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3466.4000 3930.2400 3466.5400 ;
    END
  END RES2[54]
  PIN RES2[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.7897 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.844 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3468.4400 3930.2400 3468.5800 ;
    END
  END RES2[53]
  PIN RES2[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9817 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.841 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3469.4600 3930.2400 3469.6000 ;
    END
  END RES2[52]
  PIN RES2[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.2065 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.928 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3215.4800 3930.2400 3215.6200 ;
    END
  END RES2[51]
  PIN RES2[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6941 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.403 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3216.8400 3930.2400 3216.9800 ;
    END
  END RES2[50]
  PIN RES2[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5681 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.773 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3218.5400 3930.2400 3218.6800 ;
    END
  END RES2[49]
  PIN RES2[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.0797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.331 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 3219.9000 3930.2400 3220.0400 ;
    END
  END RES2[48]
  PIN RES2[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.0777 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.284 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2965.5800 3930.2400 2965.7200 ;
    END
  END RES2[47]
  PIN RES2[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2966.9400 3930.2400 2967.0800 ;
    END
  END RES2[46]
  PIN RES2[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5037 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.451 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2968.6400 3930.2400 2968.7800 ;
    END
  END RES2[45]
  PIN RES2[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.0365 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.078 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2970.0000 3930.2400 2970.1400 ;
    END
  END RES2[44]
  PIN RES2[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2715.6800 3930.2400 2715.8200 ;
    END
  END RES2[43]
  PIN RES2[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3441 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.653 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2717.0400 3930.2400 2717.1800 ;
    END
  END RES2[42]
  PIN RES2[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6157 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.011 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2718.7400 3930.2400 2718.8800 ;
    END
  END RES2[41]
  PIN RES2[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.7949 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.907 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2720.1000 3930.2400 2720.2400 ;
    END
  END RES2[40]
  PIN RES2[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5177 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.521 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2465.7800 3930.2400 2465.9200 ;
    END
  END RES2[39]
  PIN RES2[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.2117 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.991 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2467.1400 3930.2400 2467.2800 ;
    END
  END RES2[38]
  PIN RES2[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2461 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.163 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2468.8400 3930.2400 2468.9800 ;
    END
  END RES2[37]
  PIN RES2[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.7549 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.707 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2470.2000 3930.2400 2470.3400 ;
    END
  END RES2[36]
  PIN RES2[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.1041 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.416 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2215.8800 3930.2400 2216.0200 ;
    END
  END RES2[35]
  PIN RES2[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7757 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2217.2400 3930.2400 2217.3800 ;
    END
  END RES2[34]
  PIN RES2[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6969 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.417 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2218.9400 3930.2400 2219.0800 ;
    END
  END RES2[33]
  PIN RES2[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2629 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.247 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 2220.3000 3930.2400 2220.4400 ;
    END
  END RES2[32]
  PIN RES2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.7581 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.723 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1965.9800 3930.2400 1966.1200 ;
    END
  END RES2[31]
  PIN RES2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1817 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.841 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1967.3400 3930.2400 1967.4800 ;
    END
  END RES2[30]
  PIN RES2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.5953 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.909 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1969.0400 3930.2400 1969.1800 ;
    END
  END RES2[29]
  PIN RES2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1173 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.519 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1970.4000 3930.2400 1970.5400 ;
    END
  END RES2[28]
  PIN RES2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1817 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.841 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1716.4200 3930.2400 1716.5600 ;
    END
  END RES2[27]
  PIN RES2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1717.4400 3930.2400 1717.5800 ;
    END
  END RES2[26]
  PIN RES2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7981 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.923 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1719.4800 3930.2400 1719.6200 ;
    END
  END RES2[25]
  PIN RES2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.9481 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.673 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1720.5000 3930.2400 1720.6400 ;
    END
  END RES2[24]
  PIN RES2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.769 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1466.5200 3930.2400 1466.6600 ;
    END
  END RES2[23]
  PIN RES2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2125 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.995 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1467.8800 3930.2400 1468.0200 ;
    END
  END RES2[22]
  PIN RES2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6609 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1469.5800 3930.2400 1469.7200 ;
    END
  END RES2[21]
  PIN RES2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.1441 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.653 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1470.9400 3930.2400 1471.0800 ;
    END
  END RES2[20]
  PIN RES2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3885 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.875 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1216.6200 3930.2400 1216.7600 ;
    END
  END RES2[19]
  PIN RES2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.7505 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.685 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1217.9800 3930.2400 1218.1200 ;
    END
  END RES2[18]
  PIN RES2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.8201 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.996 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1219.6800 3930.2400 1219.8200 ;
    END
  END RES2[17]
  PIN RES2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.6553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.209 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 1221.0400 3930.2400 1221.1800 ;
    END
  END RES2[16]
  PIN RES2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0497 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.181 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 966.7200 3930.2400 966.8600 ;
    END
  END RES2[15]
  PIN RES2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.8149 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.007 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 968.0800 3930.2400 968.2200 ;
    END
  END RES2[14]
  PIN RES2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.9037 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.451 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 969.7800 3930.2400 969.9200 ;
    END
  END RES2[13]
  PIN RES2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5373 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.619 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 971.1400 3930.2400 971.2800 ;
    END
  END RES2[12]
  PIN RES2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1957 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.911 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 716.8200 3930.2400 716.9600 ;
    END
  END RES2[11]
  PIN RES2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3441 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.653 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 718.1800 3930.2400 718.3200 ;
    END
  END RES2[10]
  PIN RES2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.6107 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.949 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 719.8800 3930.2400 720.0200 ;
    END
  END RES2[9]
  PIN RES2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.4393 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.129 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 721.2400 3930.2400 721.3800 ;
    END
  END RES2[8]
  PIN RES2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.4669 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.267 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 466.9200 3930.2400 467.0600 ;
    END
  END RES2[7]
  PIN RES2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.4053 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.959 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 468.2800 3930.2400 468.4200 ;
    END
  END RES2[6]
  PIN RES2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.5857 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.824 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 469.9800 3930.2400 470.1200 ;
    END
  END RES2[5]
  PIN RES2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.2997 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.431 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 471.3400 3930.2400 471.4800 ;
    END
  END RES2[4]
  PIN RES2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 217.3600 3930.2400 217.5000 ;
    END
  END RES2[3]
  PIN RES2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0497 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.181 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 218.7200 3930.2400 218.8600 ;
    END
  END RES2[2]
  PIN RES2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0221 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.043 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 220.4200 3930.2400 220.5600 ;
    END
  END RES2[1]
  PIN RES2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.1445 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.655 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 3929.6450 221.7800 3930.2400 221.9200 ;
    END
  END RES2[0]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 68.048 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 109.752 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met5  ;
    ANTENNAMAXAREACAR 71.6111 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 325.345 LAYER met5  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1791.5600 0.5950 1791.7000 ;
    END
  END CLK
  PIN SelfWriteStrobe
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 11.9432 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.1535 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1367.9600 0.8000 1368.2600 ;
    END
  END SelfWriteStrobe
  PIN SelfWriteData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5713 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.789 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 13.138 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 54.9657 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1422.3200 0.5950 1422.4600 ;
    END
  END SelfWriteData[31]
  PIN SelfWriteData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4425 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 11.8345 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 51.4424 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1425.3800 0.5950 1425.5200 ;
    END
  END SelfWriteData[30]
  PIN SelfWriteData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5069 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.467 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.4943 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 50.8606 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1416.8800 0.5950 1417.0200 ;
    END
  END SelfWriteData[29]
  PIN SelfWriteData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4425 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.2341 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 49.5596 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1406.0000 0.5950 1406.1400 ;
    END
  END SelfWriteData[28]
  PIN SelfWriteData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3781 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.823 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 9.97394 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 48.2586 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1387.3000 0.5950 1387.4400 ;
    END
  END SelfWriteData[27]
  PIN SelfWriteData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3245 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.555 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 15.8653 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 69.8101 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1403.6200 0.5950 1403.7600 ;
    END
  END SelfWriteData[26]
  PIN SelfWriteData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 25.1376 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.477 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1387.4800 0.8000 1387.7800 ;
    END
  END SelfWriteData[25]
  PIN SelfWriteData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2765 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.315 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 18.077 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 87.1192 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1400.5600 0.5950 1400.7000 ;
    END
  END SelfWriteData[24]
  PIN SelfWriteData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 14.4341 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 68.9051 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1384.2400 0.5950 1384.3800 ;
    END
  END SelfWriteData[23]
  PIN SelfWriteData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 14.0014 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 68.396 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1395.1200 0.5950 1395.2600 ;
    END
  END SelfWriteData[22]
  PIN SelfWriteData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 36.6547 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 186.253 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1384.4300 0.8000 1384.7300 ;
    END
  END SelfWriteData[21]
  PIN SelfWriteData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4701 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.283 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 14.8188 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 70.8283 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1367.9200 0.5950 1368.0600 ;
    END
  END SelfWriteData[20]
  PIN SelfWriteData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3781 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.823 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 9.97394 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 48.2586 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1392.7400 0.5950 1392.8800 ;
    END
  END SelfWriteData[19]
  PIN SelfWriteData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 26.4022 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.156 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1400.2900 0.8000 1400.5900 ;
    END
  END SelfWriteData[18]
  PIN SelfWriteData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5377 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.621 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.6188 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 51.4828 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1399.8800 0.5950 1400.0200 ;
    END
  END SelfWriteData[17]
  PIN SelfWriteData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3917 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.891 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 14.5844 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 69.3414 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1398.1800 0.5950 1398.3200 ;
    END
  END SelfWriteData[16]
  PIN SelfWriteData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9185 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.488 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 17.7982 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 81.1111 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1381.8600 0.5950 1382.0000 ;
    END
  END SelfWriteData[15]
  PIN SelfWriteData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4425 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.2341 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 49.5596 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1414.5000 0.5950 1414.6400 ;
    END
  END SelfWriteData[14]
  PIN SelfWriteData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6357 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.111 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 11.0147 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 53.4626 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1419.9400 0.5950 1420.0800 ;
    END
  END SelfWriteData[13]
  PIN SelfWriteData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4425 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.145 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 11.8345 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 51.4424 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1409.0600 0.5950 1409.2000 ;
    END
  END SelfWriteData[12]
  PIN SelfWriteData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3749 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.807 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 14.0014 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 68.396 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1411.4400 0.5950 1411.5800 ;
    END
  END SelfWriteData[11]
  PIN SelfWriteData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 12.0273 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.3798 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1403.3400 0.8000 1403.6400 ;
    END
  END SelfWriteData[10]
  PIN SelfWriteData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 39.3364 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 207.255 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1381.9900 0.8000 1382.2900 ;
    END
  END SelfWriteData[9]
  PIN SelfWriteData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 28.837 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.008 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1392.3600 0.8000 1392.6600 ;
    END
  END SelfWriteData[8]
  PIN SelfWriteData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4089 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.977 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.5311 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 49.3899 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1381.1800 0.5950 1381.3200 ;
    END
  END SelfWriteData[7]
  PIN SelfWriteData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 24.119 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.299 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1394.8000 0.8000 1395.1000 ;
    END
  END SelfWriteData[6]
  PIN SelfWriteData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3781 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.823 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 12.0414 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 50.6909 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1376.4200 0.5950 1376.5600 ;
    END
  END SelfWriteData[5]
  PIN SelfWriteData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2493 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.179 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 12.0018 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 48.6545 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1373.3600 0.5950 1373.5000 ;
    END
  END SelfWriteData[4]
  PIN SelfWriteData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5713 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.789 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.7545 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 52.1616 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1389.6800 0.5950 1389.8200 ;
    END
  END SelfWriteData[3]
  PIN SelfWriteData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 28.5145 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 148.404 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1389.3100 0.8000 1389.6100 ;
    END
  END SelfWriteData[2]
  PIN SelfWriteData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4733 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.299 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 10.3586 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 50.1818 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1383.5600 0.5950 1383.7000 ;
    END
  END SelfWriteData[1]
  PIN SelfWriteData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2629 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.247 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met1  ;
    ANTENNAMAXAREACAR 15.3828 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 68.2909 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1370.9800 0.5950 1371.1200 ;
    END
  END SelfWriteData[0]
  PIN Rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9717 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.791 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 33.7171 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 128.778 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1577.7000 0.5950 1577.8400 ;
    END
  END Rx
  PIN ComActive
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.5037 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.414 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1401.2400 0.5950 1401.3800 ;
    END
  END ComActive
  PIN ReceiveLED
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3137 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.501 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1378.4600 0.5950 1378.6000 ;
    END
  END ReceiveLED
  PIN s_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3137 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.501 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 20.5345 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 93.3016 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1324.4000 0.5950 1324.5400 ;
    END
  END s_clk
  PIN s_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5419 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.642 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 25.7187 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 106.325 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 1329.8400 0.5950 1329.9800 ;
    END
  END s_data
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2.0000 2.0000 6.0000 3928.0600 ;
        RECT 121.1800 133.5000 123.1800 3633.2600 ;
        RECT 157.0800 133.5000 159.0800 3633.2600 ;
        RECT 397.6400 82.9800 399.6400 3928.0600 ;
        RECT 638.1000 82.9800 640.1000 3928.0600 ;
        RECT 878.5600 82.9800 880.5600 3928.0600 ;
        RECT 1119.0200 82.9800 1121.0200 3928.0600 ;
        RECT 1359.4800 82.9800 1361.4800 3928.0600 ;
        RECT 1599.9400 82.9800 1601.9400 3928.0600 ;
        RECT 1840.4000 82.9800 1842.4000 3928.0600 ;
        RECT 2080.8600 82.9800 2082.8600 3928.0600 ;
        RECT 2321.3200 82.9800 2323.3200 3928.0600 ;
        RECT 2561.7800 82.9800 2563.7800 3928.0600 ;
        RECT 2802.2400 82.9800 2804.2400 3928.0600 ;
        RECT 3774.0800 1884.1200 3776.0800 2117.9600 ;
        RECT 3924.2400 2.0000 3928.2400 3928.0600 ;
        RECT 3042.7000 82.9800 3044.7000 3928.0600 ;
        RECT 3283.1600 82.9800 3285.1600 3928.0600 ;
        RECT 3523.6200 82.9800 3525.6200 3928.0600 ;
        RECT 3764.0800 82.9800 3766.0800 3928.0600 ;
        RECT 3813.9800 1882.1200 3815.9800 2117.9600 ;
        RECT 157.1800 82.9800 159.1800 119.2400 ;
        RECT 157.0800 133.2400 159.0800 135.5000 ;
        RECT 150.8400 142.9300 159.0800 144.4300 ;
        RECT 387.5800 133.2400 389.5800 144.6700 ;
        RECT 150.8400 392.7700 159.0800 394.2700 ;
        RECT 387.5800 383.0800 389.5800 394.5100 ;
        RECT 628.0400 133.2400 630.0400 144.6700 ;
        RECT 868.5000 133.2400 870.5000 144.6700 ;
        RECT 868.5000 383.0800 870.5000 394.5100 ;
        RECT 628.0400 383.0800 630.0400 394.5100 ;
        RECT 150.8400 642.6100 159.0800 644.1100 ;
        RECT 387.5800 632.9200 389.5800 644.3500 ;
        RECT 150.8400 892.4500 159.0800 893.9500 ;
        RECT 387.5800 882.7600 389.5800 894.1900 ;
        RECT 628.0400 632.9200 630.0400 644.3500 ;
        RECT 868.5000 632.9200 870.5000 644.3500 ;
        RECT 868.5000 882.7600 870.5000 894.1900 ;
        RECT 628.0400 882.7600 630.0400 894.1900 ;
        RECT 1108.9600 133.2400 1110.9600 144.6700 ;
        RECT 1349.4200 133.2400 1351.4200 144.6700 ;
        RECT 1349.4200 383.0800 1351.4200 394.5100 ;
        RECT 1108.9600 383.0800 1110.9600 394.5100 ;
        RECT 1589.8800 133.2400 1591.8800 144.6700 ;
        RECT 1830.3400 133.2400 1832.3400 144.6700 ;
        RECT 1830.3400 383.0800 1832.3400 394.5100 ;
        RECT 1589.8800 383.0800 1591.8800 394.5100 ;
        RECT 1349.4200 632.9200 1351.4200 644.3500 ;
        RECT 1108.9600 632.9200 1110.9600 644.3500 ;
        RECT 1349.4200 882.7600 1351.4200 894.1900 ;
        RECT 1108.9600 882.7600 1110.9600 894.1900 ;
        RECT 1589.8800 632.9200 1591.8800 644.3500 ;
        RECT 1830.3400 632.9200 1832.3400 644.3500 ;
        RECT 1589.8800 882.7600 1591.8800 894.1900 ;
        RECT 1830.3400 882.7600 1832.3400 894.1900 ;
        RECT 150.8400 1142.2900 159.0800 1143.7900 ;
        RECT 387.5800 1132.6000 389.5800 1144.0300 ;
        RECT 150.8400 1392.1300 159.0800 1393.6300 ;
        RECT 387.5800 1382.4400 389.5800 1393.8700 ;
        RECT 868.5000 1132.6000 870.5000 1144.0300 ;
        RECT 628.0400 1132.6000 630.0400 1144.0300 ;
        RECT 868.5000 1382.4400 870.5000 1393.8700 ;
        RECT 628.0400 1382.4400 630.0400 1393.8700 ;
        RECT 150.8400 1641.9700 159.0800 1643.4700 ;
        RECT 387.5800 1632.2800 389.5800 1643.7100 ;
        RECT 150.8400 1891.8100 159.0800 1893.3100 ;
        RECT 387.5800 1882.1200 389.5800 1893.5500 ;
        RECT 868.5000 1632.2800 870.5000 1643.7100 ;
        RECT 628.0400 1632.2800 630.0400 1643.7100 ;
        RECT 628.0400 1882.1200 630.0400 1893.5500 ;
        RECT 868.5000 1882.1200 870.5000 1893.5500 ;
        RECT 1349.4200 1132.6000 1351.4200 1144.0300 ;
        RECT 1108.9600 1132.6000 1110.9600 1144.0300 ;
        RECT 1349.4200 1382.4400 1351.4200 1393.8700 ;
        RECT 1108.9600 1382.4400 1110.9600 1393.8700 ;
        RECT 1589.8800 1132.6000 1591.8800 1144.0300 ;
        RECT 1830.3400 1132.6000 1832.3400 1144.0300 ;
        RECT 1589.8800 1382.4400 1591.8800 1393.8700 ;
        RECT 1830.3400 1382.4400 1832.3400 1393.8700 ;
        RECT 1349.4200 1632.2800 1351.4200 1643.7100 ;
        RECT 1108.9600 1632.2800 1110.9600 1643.7100 ;
        RECT 1108.9600 1882.1200 1110.9600 1893.5500 ;
        RECT 1349.4200 1882.1200 1351.4200 1893.5500 ;
        RECT 1589.8800 1632.2800 1591.8800 1643.7100 ;
        RECT 1830.3400 1632.2800 1832.3400 1643.7100 ;
        RECT 1830.3400 1882.1200 1832.3400 1893.5500 ;
        RECT 1589.8800 1882.1200 1591.8800 1893.5500 ;
        RECT 3813.9800 882.7600 3815.9800 1118.6000 ;
        RECT 3774.0800 884.7600 3776.0800 1118.6000 ;
        RECT 2070.8000 133.2400 2072.8000 144.6700 ;
        RECT 2311.2600 133.2400 2313.2600 144.6700 ;
        RECT 2311.2600 383.0800 2313.2600 394.5100 ;
        RECT 2070.8000 383.0800 2072.8000 394.5100 ;
        RECT 2551.7200 133.2400 2553.7200 144.6700 ;
        RECT 2792.1800 133.2400 2794.1800 144.6700 ;
        RECT 2792.1800 383.0800 2794.1800 394.5100 ;
        RECT 2551.7200 383.0800 2553.7200 394.5100 ;
        RECT 2311.2600 632.9200 2313.2600 644.3500 ;
        RECT 2070.8000 632.9200 2072.8000 644.3500 ;
        RECT 2311.2600 882.7600 2313.2600 894.1900 ;
        RECT 2070.8000 882.7600 2072.8000 894.1900 ;
        RECT 2792.1800 632.9200 2794.1800 644.3500 ;
        RECT 2551.7200 632.9200 2553.7200 644.3500 ;
        RECT 2792.1800 882.7600 2794.1800 894.1900 ;
        RECT 2551.7200 882.7600 2553.7200 894.1900 ;
        RECT 3813.9800 383.0800 3815.9800 618.9200 ;
        RECT 3774.0800 385.0800 3776.0800 618.9200 ;
        RECT 3032.6400 133.2400 3034.6400 144.6700 ;
        RECT 3273.1000 133.2400 3275.1000 144.6700 ;
        RECT 3032.6400 383.0800 3034.6400 394.5100 ;
        RECT 3273.1000 383.0800 3275.1000 394.5100 ;
        RECT 3813.9800 133.2400 3815.9800 369.0800 ;
        RECT 3774.0800 135.2400 3776.0800 369.0800 ;
        RECT 3537.6800 133.2400 3539.6800 144.6700 ;
        RECT 3513.5600 133.2400 3515.5600 144.6700 ;
        RECT 3807.7400 142.6700 3815.9800 144.1700 ;
        RECT 3513.5600 383.0800 3515.5600 394.5100 ;
        RECT 3754.0200 383.0800 3756.0200 394.5100 ;
        RECT 3807.7400 392.5100 3815.9800 394.0100 ;
        RECT 3273.1000 632.9200 3275.1000 644.3500 ;
        RECT 3032.6400 632.9200 3034.6400 644.3500 ;
        RECT 3273.1000 882.7600 3275.1000 894.1900 ;
        RECT 3032.6400 882.7600 3034.6400 894.1900 ;
        RECT 3774.0800 634.9200 3776.0800 868.7600 ;
        RECT 3813.9800 632.9200 3815.9800 868.7600 ;
        RECT 3513.5600 632.9200 3515.5600 644.3500 ;
        RECT 3754.0200 632.9200 3756.0200 644.3500 ;
        RECT 3807.7400 642.3500 3815.9800 643.8500 ;
        RECT 3513.5600 882.7600 3515.5600 894.1900 ;
        RECT 3754.0200 882.7600 3756.0200 894.1900 ;
        RECT 3807.7400 892.1900 3815.9800 893.6900 ;
        RECT 2311.2600 1132.6000 2313.2600 1144.0300 ;
        RECT 2070.8000 1132.6000 2072.8000 1144.0300 ;
        RECT 2311.2600 1382.4400 2313.2600 1393.8700 ;
        RECT 2070.8000 1382.4400 2072.8000 1393.8700 ;
        RECT 2792.1800 1132.6000 2794.1800 1144.0300 ;
        RECT 2551.7200 1132.6000 2553.7200 1144.0300 ;
        RECT 2792.1800 1382.4400 2794.1800 1393.8700 ;
        RECT 2551.7200 1382.4400 2553.7200 1393.8700 ;
        RECT 2311.2600 1632.2800 2313.2600 1643.7100 ;
        RECT 2070.8000 1632.2800 2072.8000 1643.7100 ;
        RECT 2311.2600 1882.1200 2313.2600 1893.5500 ;
        RECT 2070.8000 1882.1200 2072.8000 1893.5500 ;
        RECT 2792.1800 1632.2800 2794.1800 1643.7100 ;
        RECT 2551.7200 1632.2800 2553.7200 1643.7100 ;
        RECT 2792.1800 1882.1200 2794.1800 1893.5500 ;
        RECT 2551.7200 1882.1200 2553.7200 1893.5500 ;
        RECT 3813.9800 1382.4400 3815.9800 1618.2800 ;
        RECT 3774.0800 1384.4400 3776.0800 1618.2800 ;
        RECT 3273.1000 1132.6000 3275.1000 1144.0300 ;
        RECT 3032.6400 1132.6000 3034.6400 1144.0300 ;
        RECT 3273.1000 1382.4400 3275.1000 1393.8700 ;
        RECT 3032.6400 1382.4400 3034.6400 1393.8700 ;
        RECT 3774.0800 1134.6000 3776.0800 1368.4400 ;
        RECT 3813.9800 1132.6000 3815.9800 1368.4400 ;
        RECT 3513.5600 1132.6000 3515.5600 1144.0300 ;
        RECT 3754.0200 1132.6000 3756.0200 1144.0300 ;
        RECT 3807.7400 1142.0300 3815.9800 1143.5300 ;
        RECT 3513.5600 1382.4400 3515.5600 1393.8700 ;
        RECT 3754.0200 1382.4400 3756.0200 1393.8700 ;
        RECT 3807.7400 1391.8700 3815.9800 1393.3700 ;
        RECT 3273.1000 1632.2800 3275.1000 1643.7100 ;
        RECT 3032.6400 1632.2800 3034.6400 1643.7100 ;
        RECT 3273.1000 1882.1200 3275.1000 1893.5500 ;
        RECT 3032.6400 1882.1200 3034.6400 1893.5500 ;
        RECT 3774.0800 1634.2800 3776.0800 1868.1200 ;
        RECT 3813.9800 1632.2800 3815.9800 1868.1200 ;
        RECT 3513.5600 1632.2800 3515.5600 1643.7100 ;
        RECT 3754.0200 1632.2800 3756.0200 1643.7100 ;
        RECT 3807.7400 1641.7100 3815.9800 1643.2100 ;
        RECT 3513.5600 1882.1200 3515.5600 1893.5500 ;
        RECT 3754.0200 1882.1200 3756.0200 1893.5500 ;
        RECT 3807.7400 1891.5500 3815.9800 1893.0500 ;
        RECT 150.8400 2141.6500 159.0800 2143.1500 ;
        RECT 387.5800 2131.9600 389.5800 2143.3900 ;
        RECT 150.8400 2391.4900 159.0800 2392.9900 ;
        RECT 387.5800 2381.8000 389.5800 2393.2300 ;
        RECT 868.5000 2131.9600 870.5000 2143.3900 ;
        RECT 628.0400 2131.9600 630.0400 2143.3900 ;
        RECT 868.5000 2381.8000 870.5000 2393.2300 ;
        RECT 628.0400 2381.8000 630.0400 2393.2300 ;
        RECT 150.8400 2641.3300 159.0800 2642.8300 ;
        RECT 387.5800 2631.6400 389.5800 2643.0700 ;
        RECT 150.8400 2891.1700 159.0800 2892.6700 ;
        RECT 387.5800 2881.4800 389.5800 2892.9100 ;
        RECT 868.5000 2631.6400 870.5000 2643.0700 ;
        RECT 628.0400 2631.6400 630.0400 2643.0700 ;
        RECT 868.5000 2881.4800 870.5000 2892.9100 ;
        RECT 628.0400 2881.4800 630.0400 2892.9100 ;
        RECT 1349.4200 2131.9600 1351.4200 2143.3900 ;
        RECT 1108.9600 2131.9600 1110.9600 2143.3900 ;
        RECT 1349.4200 2381.8000 1351.4200 2393.2300 ;
        RECT 1108.9600 2381.8000 1110.9600 2393.2300 ;
        RECT 1589.8800 2131.9600 1591.8800 2143.3900 ;
        RECT 1830.3400 2131.9600 1832.3400 2143.3900 ;
        RECT 1589.8800 2381.8000 1591.8800 2393.2300 ;
        RECT 1830.3400 2381.8000 1832.3400 2393.2300 ;
        RECT 1349.4200 2631.6400 1351.4200 2643.0700 ;
        RECT 1108.9600 2631.6400 1110.9600 2643.0700 ;
        RECT 1349.4200 2881.4800 1351.4200 2892.9100 ;
        RECT 1108.9600 2881.4800 1110.9600 2892.9100 ;
        RECT 1589.8800 2631.6400 1591.8800 2643.0700 ;
        RECT 1830.3400 2631.6400 1832.3400 2643.0700 ;
        RECT 1589.8800 2881.4800 1591.8800 2892.9100 ;
        RECT 1830.3400 2881.4800 1832.3400 2892.9100 ;
        RECT 150.8400 3141.0100 159.0800 3142.5100 ;
        RECT 387.5800 3131.3200 389.5800 3142.7500 ;
        RECT 150.8400 3390.8500 159.0800 3392.3500 ;
        RECT 387.5800 3381.1600 389.5800 3392.5900 ;
        RECT 628.0400 3131.3200 630.0400 3142.7500 ;
        RECT 868.5000 3131.3200 870.5000 3142.7500 ;
        RECT 628.0400 3381.1600 630.0400 3392.5900 ;
        RECT 868.5000 3381.1600 870.5000 3392.5900 ;
        RECT 121.1800 3631.2600 123.1800 3928.0600 ;
        RECT 157.0800 3631.2600 159.0800 3928.0600 ;
        RECT 150.8400 3640.6900 159.0800 3642.1900 ;
        RECT 387.5800 3631.0000 389.5800 3642.4300 ;
        RECT 397.6400 3882.8400 399.6400 3928.0600 ;
        RECT 868.5000 3631.0000 870.5000 3642.4300 ;
        RECT 628.0400 3631.0000 630.0400 3642.4300 ;
        RECT 638.1000 3882.8400 640.1000 3928.0600 ;
        RECT 878.5600 3882.8400 880.5600 3928.0600 ;
        RECT 1349.4200 3131.3200 1351.4200 3142.7500 ;
        RECT 1108.9600 3131.3200 1110.9600 3142.7500 ;
        RECT 1349.4200 3381.1600 1351.4200 3392.5900 ;
        RECT 1108.9600 3381.1600 1110.9600 3392.5900 ;
        RECT 1589.8800 3131.3200 1591.8800 3142.7500 ;
        RECT 1830.3400 3131.3200 1832.3400 3142.7500 ;
        RECT 1589.8800 3381.1600 1591.8800 3392.5900 ;
        RECT 1830.3400 3381.1600 1832.3400 3392.5900 ;
        RECT 1108.9600 3631.0000 1110.9600 3642.4300 ;
        RECT 1349.4200 3631.0000 1351.4200 3642.4300 ;
        RECT 1119.0200 3882.8400 1121.0200 3928.0600 ;
        RECT 1359.4800 3882.8400 1361.4800 3928.0600 ;
        RECT 1830.3400 3631.0000 1832.3400 3642.4300 ;
        RECT 1589.8800 3631.0000 1591.8800 3642.4300 ;
        RECT 1599.9400 3882.8400 1601.9400 3928.0600 ;
        RECT 1840.4000 3882.8400 1842.4000 3928.0600 ;
        RECT 3813.9800 2881.4800 3815.9800 3117.3200 ;
        RECT 3774.0800 2883.4800 3776.0800 3117.3200 ;
        RECT 2311.2600 2131.9600 2313.2600 2143.3900 ;
        RECT 2070.8000 2131.9600 2072.8000 2143.3900 ;
        RECT 2311.2600 2381.8000 2313.2600 2393.2300 ;
        RECT 2070.8000 2381.8000 2072.8000 2393.2300 ;
        RECT 2792.1800 2131.9600 2794.1800 2143.3900 ;
        RECT 2551.7200 2131.9600 2553.7200 2143.3900 ;
        RECT 2792.1800 2381.8000 2794.1800 2393.2300 ;
        RECT 2551.7200 2381.8000 2553.7200 2393.2300 ;
        RECT 2311.2600 2631.6400 2313.2600 2643.0700 ;
        RECT 2070.8000 2631.6400 2072.8000 2643.0700 ;
        RECT 2311.2600 2881.4800 2313.2600 2892.9100 ;
        RECT 2070.8000 2881.4800 2072.8000 2892.9100 ;
        RECT 2792.1800 2631.6400 2794.1800 2643.0700 ;
        RECT 2551.7200 2631.6400 2553.7200 2643.0700 ;
        RECT 2792.1800 2881.4800 2794.1800 2892.9100 ;
        RECT 2551.7200 2881.4800 2553.7200 2892.9100 ;
        RECT 3813.9800 2381.8000 3815.9800 2617.6400 ;
        RECT 3774.0800 2383.8000 3776.0800 2617.6400 ;
        RECT 3273.1000 2131.9600 3275.1000 2143.3900 ;
        RECT 3032.6400 2131.9600 3034.6400 2143.3900 ;
        RECT 3273.1000 2381.8000 3275.1000 2393.2300 ;
        RECT 3032.6400 2381.8000 3034.6400 2393.2300 ;
        RECT 3774.0800 2133.9600 3776.0800 2367.8000 ;
        RECT 3813.9800 2131.9600 3815.9800 2367.8000 ;
        RECT 3513.5600 2131.9600 3515.5600 2143.3900 ;
        RECT 3754.0200 2131.9600 3756.0200 2143.3900 ;
        RECT 3807.7400 2141.3900 3815.9800 2142.8900 ;
        RECT 3513.5600 2381.8000 3515.5600 2393.2300 ;
        RECT 3754.0200 2381.8000 3756.0200 2393.2300 ;
        RECT 3807.7400 2391.2300 3815.9800 2392.7300 ;
        RECT 3273.1000 2631.6400 3275.1000 2643.0700 ;
        RECT 3032.6400 2631.6400 3034.6400 2643.0700 ;
        RECT 3273.1000 2881.4800 3275.1000 2892.9100 ;
        RECT 3032.6400 2881.4800 3034.6400 2892.9100 ;
        RECT 3774.0800 2633.6400 3776.0800 2867.4800 ;
        RECT 3813.9800 2631.6400 3815.9800 2867.4800 ;
        RECT 3513.5600 2631.6400 3515.5600 2643.0700 ;
        RECT 3754.0200 2631.6400 3756.0200 2643.0700 ;
        RECT 3807.7400 2641.0700 3815.9800 2642.5700 ;
        RECT 3513.5600 2881.4800 3515.5600 2892.9100 ;
        RECT 3754.0200 2881.4800 3756.0200 2892.9100 ;
        RECT 3807.7400 2890.9100 3815.9800 2892.4100 ;
        RECT 2311.2600 3131.3200 2313.2600 3142.7500 ;
        RECT 2070.8000 3131.3200 2072.8000 3142.7500 ;
        RECT 2311.2600 3381.1600 2313.2600 3392.5900 ;
        RECT 2070.8000 3381.1600 2072.8000 3392.5900 ;
        RECT 2792.1800 3131.3200 2794.1800 3142.7500 ;
        RECT 2551.7200 3131.3200 2553.7200 3142.7500 ;
        RECT 2792.1800 3381.1600 2794.1800 3392.5900 ;
        RECT 2551.7200 3381.1600 2553.7200 3392.5900 ;
        RECT 2070.8000 3631.0000 2072.8000 3642.4300 ;
        RECT 2311.2600 3631.0000 2313.2600 3642.4300 ;
        RECT 2080.8600 3882.8400 2082.8600 3928.0600 ;
        RECT 2321.3200 3882.8400 2323.3200 3928.0600 ;
        RECT 2551.7200 3631.0000 2553.7200 3642.4300 ;
        RECT 2561.7800 3882.8400 2563.7800 3928.0600 ;
        RECT 2802.2400 3882.8400 2804.2400 3928.0600 ;
        RECT 3813.9800 3381.1600 3815.9800 3617.0000 ;
        RECT 3774.0800 3383.1600 3776.0800 3617.0000 ;
        RECT 3273.1000 3131.3200 3275.1000 3142.7500 ;
        RECT 3032.6400 3131.3200 3034.6400 3142.7500 ;
        RECT 3273.1000 3381.1600 3275.1000 3392.5900 ;
        RECT 3032.6400 3381.1600 3034.6400 3392.5900 ;
        RECT 3774.0800 3133.3200 3776.0800 3367.1600 ;
        RECT 3813.9800 3131.3200 3815.9800 3367.1600 ;
        RECT 3513.5600 3131.3200 3515.5600 3142.7500 ;
        RECT 3754.0200 3131.3200 3756.0200 3142.7500 ;
        RECT 3807.7400 3140.7500 3815.9800 3142.2500 ;
        RECT 3513.5600 3381.1600 3515.5600 3392.5900 ;
        RECT 3754.0200 3381.1600 3756.0200 3392.5900 ;
        RECT 3807.7400 3390.5900 3815.9800 3392.0900 ;
        RECT 3032.6400 3631.0000 3034.6400 3642.4300 ;
        RECT 3273.1000 3631.0000 3275.1000 3642.4300 ;
        RECT 3042.7000 3882.8400 3044.7000 3928.0600 ;
        RECT 3283.1600 3882.8400 3285.1600 3928.0600 ;
        RECT 3813.9800 3631.0000 3815.9800 3866.8400 ;
        RECT 3774.0800 3633.0000 3776.0800 3866.8400 ;
        RECT 3513.5600 3631.0000 3515.5600 3642.4300 ;
        RECT 3754.0200 3631.0000 3756.0200 3642.4300 ;
        RECT 3807.7400 3640.4300 3815.9800 3641.9300 ;
        RECT 3523.6200 3882.8400 3525.6200 3928.0600 ;
        RECT 3764.0800 3882.8400 3766.0800 3928.0600 ;
        RECT 150.0900 142.9300 151.5900 144.4300 ;
        RECT 387.5800 143.1700 389.5800 145.6700 ;
        RECT 150.0900 392.7700 151.5900 394.2700 ;
        RECT 387.5800 393.0100 389.5800 395.5100 ;
        RECT 628.0400 143.1700 630.0400 145.6700 ;
        RECT 868.5000 143.1700 870.5000 145.6700 ;
        RECT 628.0400 393.0100 630.0400 395.5100 ;
        RECT 868.5000 393.0100 870.5000 395.5100 ;
        RECT 150.0900 642.6100 151.5900 644.1100 ;
        RECT 387.5800 642.8500 389.5800 645.3500 ;
        RECT 150.0900 892.4500 151.5900 893.9500 ;
        RECT 387.5800 892.6900 389.5800 895.1900 ;
        RECT 628.0400 642.8500 630.0400 645.3500 ;
        RECT 868.5000 642.8500 870.5000 645.3500 ;
        RECT 628.0400 892.6900 630.0400 895.1900 ;
        RECT 868.5000 892.6900 870.5000 895.1900 ;
        RECT 1108.9600 143.1700 1110.9600 145.6700 ;
        RECT 1349.4200 143.1700 1351.4200 145.6700 ;
        RECT 1108.9600 393.0100 1110.9600 395.5100 ;
        RECT 1349.4200 393.0100 1351.4200 395.5100 ;
        RECT 1589.8800 143.1700 1591.8800 145.6700 ;
        RECT 1830.3400 143.1700 1832.3400 145.6700 ;
        RECT 1589.8800 393.0100 1591.8800 395.5100 ;
        RECT 1830.3400 393.0100 1832.3400 395.5100 ;
        RECT 1108.9600 642.8500 1110.9600 645.3500 ;
        RECT 1349.4200 642.8500 1351.4200 645.3500 ;
        RECT 1108.9600 892.6900 1110.9600 895.1900 ;
        RECT 1349.4200 892.6900 1351.4200 895.1900 ;
        RECT 1589.8800 642.8500 1591.8800 645.3500 ;
        RECT 1830.3400 642.8500 1832.3400 645.3500 ;
        RECT 1589.8800 892.6900 1591.8800 895.1900 ;
        RECT 1830.3400 892.6900 1832.3400 895.1900 ;
        RECT 150.0900 1142.2900 151.5900 1143.7900 ;
        RECT 387.5800 1142.5300 389.5800 1145.0300 ;
        RECT 150.0900 1392.1300 151.5900 1393.6300 ;
        RECT 387.5800 1392.3700 389.5800 1394.8700 ;
        RECT 628.0400 1142.5300 630.0400 1145.0300 ;
        RECT 868.5000 1142.5300 870.5000 1145.0300 ;
        RECT 628.0400 1392.3700 630.0400 1394.8700 ;
        RECT 868.5000 1392.3700 870.5000 1394.8700 ;
        RECT 150.0900 1641.9700 151.5900 1643.4700 ;
        RECT 387.5800 1642.2100 389.5800 1644.7100 ;
        RECT 150.0900 1891.8100 151.5900 1893.3100 ;
        RECT 387.5800 1892.0500 389.5800 1894.5500 ;
        RECT 628.0400 1642.2100 630.0400 1644.7100 ;
        RECT 868.5000 1642.2100 870.5000 1644.7100 ;
        RECT 628.0400 1892.0500 630.0400 1894.5500 ;
        RECT 868.5000 1892.0500 870.5000 1894.5500 ;
        RECT 1108.9600 1142.5300 1110.9600 1145.0300 ;
        RECT 1349.4200 1142.5300 1351.4200 1145.0300 ;
        RECT 1108.9600 1392.3700 1110.9600 1394.8700 ;
        RECT 1349.4200 1392.3700 1351.4200 1394.8700 ;
        RECT 1589.8800 1142.5300 1591.8800 1145.0300 ;
        RECT 1830.3400 1142.5300 1832.3400 1145.0300 ;
        RECT 1589.8800 1392.3700 1591.8800 1394.8700 ;
        RECT 1830.3400 1392.3700 1832.3400 1394.8700 ;
        RECT 1108.9600 1642.2100 1110.9600 1644.7100 ;
        RECT 1349.4200 1642.2100 1351.4200 1644.7100 ;
        RECT 1108.9600 1892.0500 1110.9600 1894.5500 ;
        RECT 1349.4200 1892.0500 1351.4200 1894.5500 ;
        RECT 1589.8800 1642.2100 1591.8800 1644.7100 ;
        RECT 1830.3400 1642.2100 1832.3400 1644.7100 ;
        RECT 1589.8800 1892.0500 1591.8800 1894.5500 ;
        RECT 1830.3400 1892.0500 1832.3400 1894.5500 ;
        RECT 2070.8000 143.1700 2072.8000 145.6700 ;
        RECT 2311.2600 143.1700 2313.2600 145.6700 ;
        RECT 2070.8000 393.0100 2072.8000 395.5100 ;
        RECT 2311.2600 393.0100 2313.2600 395.5100 ;
        RECT 2551.7200 143.1700 2553.7200 145.6700 ;
        RECT 2792.1800 143.1700 2794.1800 145.6700 ;
        RECT 2551.7200 393.0100 2553.7200 395.5100 ;
        RECT 2792.1800 393.0100 2794.1800 395.5100 ;
        RECT 2070.8000 642.8500 2072.8000 645.3500 ;
        RECT 2311.2600 642.8500 2313.2600 645.3500 ;
        RECT 2070.8000 892.6900 2072.8000 895.1900 ;
        RECT 2311.2600 892.6900 2313.2600 895.1900 ;
        RECT 2551.7200 642.8500 2553.7200 645.3500 ;
        RECT 2792.1800 642.8500 2794.1800 645.3500 ;
        RECT 2551.7200 892.6900 2553.7200 895.1900 ;
        RECT 2792.1800 892.6900 2794.1800 895.1900 ;
        RECT 3032.6400 143.1700 3034.6400 145.6700 ;
        RECT 3273.1000 143.1700 3275.1000 145.6700 ;
        RECT 3032.6400 393.0100 3034.6400 395.5100 ;
        RECT 3273.1000 393.0100 3275.1000 395.5100 ;
        RECT 3513.5600 143.1700 3515.5600 145.6700 ;
        RECT 3537.6800 143.1700 3539.6800 145.6700 ;
        RECT 3806.9900 142.6700 3808.4900 144.1700 ;
        RECT 3513.5600 393.0100 3515.5600 395.5100 ;
        RECT 3806.9900 392.5100 3808.4900 394.0100 ;
        RECT 3754.0200 393.0100 3756.0200 395.5100 ;
        RECT 3032.6400 642.8500 3034.6400 645.3500 ;
        RECT 3273.1000 642.8500 3275.1000 645.3500 ;
        RECT 3032.6400 892.6900 3034.6400 895.1900 ;
        RECT 3273.1000 892.6900 3275.1000 895.1900 ;
        RECT 3513.5600 642.8500 3515.5600 645.3500 ;
        RECT 3806.9900 642.3500 3808.4900 643.8500 ;
        RECT 3754.0200 642.8500 3756.0200 645.3500 ;
        RECT 3513.5600 892.6900 3515.5600 895.1900 ;
        RECT 3806.9900 892.1900 3808.4900 893.6900 ;
        RECT 3754.0200 892.6900 3756.0200 895.1900 ;
        RECT 2070.8000 1142.5300 2072.8000 1145.0300 ;
        RECT 2311.2600 1142.5300 2313.2600 1145.0300 ;
        RECT 2070.8000 1392.3700 2072.8000 1394.8700 ;
        RECT 2311.2600 1392.3700 2313.2600 1394.8700 ;
        RECT 2551.7200 1142.5300 2553.7200 1145.0300 ;
        RECT 2792.1800 1142.5300 2794.1800 1145.0300 ;
        RECT 2551.7200 1392.3700 2553.7200 1394.8700 ;
        RECT 2792.1800 1392.3700 2794.1800 1394.8700 ;
        RECT 2070.8000 1642.2100 2072.8000 1644.7100 ;
        RECT 2311.2600 1642.2100 2313.2600 1644.7100 ;
        RECT 2070.8000 1892.0500 2072.8000 1894.5500 ;
        RECT 2311.2600 1892.0500 2313.2600 1894.5500 ;
        RECT 2551.7200 1642.2100 2553.7200 1644.7100 ;
        RECT 2792.1800 1642.2100 2794.1800 1644.7100 ;
        RECT 2551.7200 1892.0500 2553.7200 1894.5500 ;
        RECT 2792.1800 1892.0500 2794.1800 1894.5500 ;
        RECT 3032.6400 1142.5300 3034.6400 1145.0300 ;
        RECT 3273.1000 1142.5300 3275.1000 1145.0300 ;
        RECT 3032.6400 1392.3700 3034.6400 1394.8700 ;
        RECT 3273.1000 1392.3700 3275.1000 1394.8700 ;
        RECT 3513.5600 1142.5300 3515.5600 1145.0300 ;
        RECT 3806.9900 1142.0300 3808.4900 1143.5300 ;
        RECT 3754.0200 1142.5300 3756.0200 1145.0300 ;
        RECT 3513.5600 1392.3700 3515.5600 1394.8700 ;
        RECT 3806.9900 1391.8700 3808.4900 1393.3700 ;
        RECT 3754.0200 1392.3700 3756.0200 1394.8700 ;
        RECT 3032.6400 1642.2100 3034.6400 1644.7100 ;
        RECT 3273.1000 1642.2100 3275.1000 1644.7100 ;
        RECT 3032.6400 1892.0500 3034.6400 1894.5500 ;
        RECT 3273.1000 1892.0500 3275.1000 1894.5500 ;
        RECT 3513.5600 1642.2100 3515.5600 1644.7100 ;
        RECT 3806.9900 1641.7100 3808.4900 1643.2100 ;
        RECT 3754.0200 1642.2100 3756.0200 1644.7100 ;
        RECT 3513.5600 1892.0500 3515.5600 1894.5500 ;
        RECT 3806.9900 1891.5500 3808.4900 1893.0500 ;
        RECT 3754.0200 1892.0500 3756.0200 1894.5500 ;
        RECT 150.0900 2141.6500 151.5900 2143.1500 ;
        RECT 387.5800 2141.8900 389.5800 2144.3900 ;
        RECT 150.0900 2391.4900 151.5900 2392.9900 ;
        RECT 387.5800 2391.7300 389.5800 2394.2300 ;
        RECT 628.0400 2141.8900 630.0400 2144.3900 ;
        RECT 868.5000 2141.8900 870.5000 2144.3900 ;
        RECT 628.0400 2391.7300 630.0400 2394.2300 ;
        RECT 868.5000 2391.7300 870.5000 2394.2300 ;
        RECT 150.0900 2641.3300 151.5900 2642.8300 ;
        RECT 387.5800 2641.5700 389.5800 2644.0700 ;
        RECT 150.0900 2891.1700 151.5900 2892.6700 ;
        RECT 387.5800 2891.4100 389.5800 2893.9100 ;
        RECT 628.0400 2641.5700 630.0400 2644.0700 ;
        RECT 868.5000 2641.5700 870.5000 2644.0700 ;
        RECT 628.0400 2891.4100 630.0400 2893.9100 ;
        RECT 868.5000 2891.4100 870.5000 2893.9100 ;
        RECT 1108.9600 2141.8900 1110.9600 2144.3900 ;
        RECT 1349.4200 2141.8900 1351.4200 2144.3900 ;
        RECT 1108.9600 2391.7300 1110.9600 2394.2300 ;
        RECT 1349.4200 2391.7300 1351.4200 2394.2300 ;
        RECT 1589.8800 2141.8900 1591.8800 2144.3900 ;
        RECT 1830.3400 2141.8900 1832.3400 2144.3900 ;
        RECT 1589.8800 2391.7300 1591.8800 2394.2300 ;
        RECT 1830.3400 2391.7300 1832.3400 2394.2300 ;
        RECT 1108.9600 2641.5700 1110.9600 2644.0700 ;
        RECT 1349.4200 2641.5700 1351.4200 2644.0700 ;
        RECT 1108.9600 2891.4100 1110.9600 2893.9100 ;
        RECT 1349.4200 2891.4100 1351.4200 2893.9100 ;
        RECT 1589.8800 2641.5700 1591.8800 2644.0700 ;
        RECT 1830.3400 2641.5700 1832.3400 2644.0700 ;
        RECT 1589.8800 2891.4100 1591.8800 2893.9100 ;
        RECT 1830.3400 2891.4100 1832.3400 2893.9100 ;
        RECT 150.0900 3141.0100 151.5900 3142.5100 ;
        RECT 387.5800 3141.2500 389.5800 3143.7500 ;
        RECT 150.0900 3390.8500 151.5900 3392.3500 ;
        RECT 387.5800 3391.0900 389.5800 3393.5900 ;
        RECT 628.0400 3141.2500 630.0400 3143.7500 ;
        RECT 868.5000 3141.2500 870.5000 3143.7500 ;
        RECT 628.0400 3391.0900 630.0400 3393.5900 ;
        RECT 868.5000 3391.0900 870.5000 3393.5900 ;
        RECT 150.0900 3640.6900 151.5900 3642.1900 ;
        RECT 387.5800 3640.9300 389.5800 3643.4300 ;
        RECT 628.0400 3640.9300 630.0400 3643.4300 ;
        RECT 868.5000 3640.9300 870.5000 3643.4300 ;
        RECT 1108.9600 3141.2500 1110.9600 3143.7500 ;
        RECT 1349.4200 3141.2500 1351.4200 3143.7500 ;
        RECT 1108.9600 3391.0900 1110.9600 3393.5900 ;
        RECT 1349.4200 3391.0900 1351.4200 3393.5900 ;
        RECT 1589.8800 3141.2500 1591.8800 3143.7500 ;
        RECT 1830.3400 3141.2500 1832.3400 3143.7500 ;
        RECT 1589.8800 3391.0900 1591.8800 3393.5900 ;
        RECT 1830.3400 3391.0900 1832.3400 3393.5900 ;
        RECT 1108.9600 3640.9300 1110.9600 3643.4300 ;
        RECT 1349.4200 3640.9300 1351.4200 3643.4300 ;
        RECT 1589.8800 3640.9300 1591.8800 3643.4300 ;
        RECT 1830.3400 3640.9300 1832.3400 3643.4300 ;
        RECT 2070.8000 2141.8900 2072.8000 2144.3900 ;
        RECT 2311.2600 2141.8900 2313.2600 2144.3900 ;
        RECT 2070.8000 2391.7300 2072.8000 2394.2300 ;
        RECT 2311.2600 2391.7300 2313.2600 2394.2300 ;
        RECT 2551.7200 2141.8900 2553.7200 2144.3900 ;
        RECT 2792.1800 2141.8900 2794.1800 2144.3900 ;
        RECT 2551.7200 2391.7300 2553.7200 2394.2300 ;
        RECT 2792.1800 2391.7300 2794.1800 2394.2300 ;
        RECT 2070.8000 2641.5700 2072.8000 2644.0700 ;
        RECT 2311.2600 2641.5700 2313.2600 2644.0700 ;
        RECT 2070.8000 2891.4100 2072.8000 2893.9100 ;
        RECT 2311.2600 2891.4100 2313.2600 2893.9100 ;
        RECT 2551.7200 2641.5700 2553.7200 2644.0700 ;
        RECT 2792.1800 2641.5700 2794.1800 2644.0700 ;
        RECT 2551.7200 2891.4100 2553.7200 2893.9100 ;
        RECT 2792.1800 2891.4100 2794.1800 2893.9100 ;
        RECT 3032.6400 2141.8900 3034.6400 2144.3900 ;
        RECT 3273.1000 2141.8900 3275.1000 2144.3900 ;
        RECT 3032.6400 2391.7300 3034.6400 2394.2300 ;
        RECT 3273.1000 2391.7300 3275.1000 2394.2300 ;
        RECT 3513.5600 2141.8900 3515.5600 2144.3900 ;
        RECT 3806.9900 2141.3900 3808.4900 2142.8900 ;
        RECT 3754.0200 2141.8900 3756.0200 2144.3900 ;
        RECT 3513.5600 2391.7300 3515.5600 2394.2300 ;
        RECT 3806.9900 2391.2300 3808.4900 2392.7300 ;
        RECT 3754.0200 2391.7300 3756.0200 2394.2300 ;
        RECT 3774.0800 2367.4950 3776.0800 2367.8250 ;
        RECT 3813.9800 2367.4950 3815.9800 2367.8250 ;
        RECT 3032.6400 2641.5700 3034.6400 2644.0700 ;
        RECT 3273.1000 2641.5700 3275.1000 2644.0700 ;
        RECT 3032.6400 2891.4100 3034.6400 2893.9100 ;
        RECT 3273.1000 2891.4100 3275.1000 2893.9100 ;
        RECT 3513.5600 2641.5700 3515.5600 2644.0700 ;
        RECT 3806.9900 2641.0700 3808.4900 2642.5700 ;
        RECT 3754.0200 2641.5700 3756.0200 2644.0700 ;
        RECT 3513.5600 2891.4100 3515.5600 2893.9100 ;
        RECT 3806.9900 2890.9100 3808.4900 2892.4100 ;
        RECT 3754.0200 2891.4100 3756.0200 2893.9100 ;
        RECT 2070.8000 3141.2500 2072.8000 3143.7500 ;
        RECT 2311.2600 3141.2500 2313.2600 3143.7500 ;
        RECT 2070.8000 3391.0900 2072.8000 3393.5900 ;
        RECT 2311.2600 3391.0900 2313.2600 3393.5900 ;
        RECT 2551.7200 3141.2500 2553.7200 3143.7500 ;
        RECT 2792.1800 3141.2500 2794.1800 3143.7500 ;
        RECT 2551.7200 3391.0900 2553.7200 3393.5900 ;
        RECT 2792.1800 3391.0900 2794.1800 3393.5900 ;
        RECT 2070.8000 3640.9300 2072.8000 3643.4300 ;
        RECT 2311.2600 3640.9300 2313.2600 3643.4300 ;
        RECT 2551.7200 3640.9300 2553.7200 3643.4300 ;
        RECT 3032.6400 3141.2500 3034.6400 3143.7500 ;
        RECT 3273.1000 3141.2500 3275.1000 3143.7500 ;
        RECT 3032.6400 3391.0900 3034.6400 3393.5900 ;
        RECT 3273.1000 3391.0900 3275.1000 3393.5900 ;
        RECT 3513.5600 3141.2500 3515.5600 3143.7500 ;
        RECT 3806.9900 3140.7500 3808.4900 3142.2500 ;
        RECT 3754.0200 3141.2500 3756.0200 3143.7500 ;
        RECT 3513.5600 3391.0900 3515.5600 3393.5900 ;
        RECT 3806.9900 3390.5900 3808.4900 3392.0900 ;
        RECT 3754.0200 3391.0900 3756.0200 3393.5900 ;
        RECT 3032.6400 3640.9300 3034.6400 3643.4300 ;
        RECT 3273.1000 3640.9300 3275.1000 3643.4300 ;
        RECT 3513.5600 3640.9300 3515.5600 3643.4300 ;
        RECT 3806.9900 3640.4300 3808.4900 3641.9300 ;
        RECT 3754.0200 3640.9300 3756.0200 3643.4300 ;
        RECT 388.0800 91.0500 390.0800 93.0500 ;
        RECT 628.5400 91.0500 630.5400 93.0500 ;
        RECT 869.0000 91.0500 871.0000 93.0500 ;
        RECT 1109.4600 91.0500 1111.4600 93.0500 ;
        RECT 1349.9200 91.0500 1351.9200 93.0500 ;
        RECT 1590.3800 91.0500 1592.3800 93.0500 ;
        RECT 1830.8400 91.0500 1832.8400 93.0500 ;
        RECT 2071.3000 91.0500 2073.3000 93.0500 ;
        RECT 2311.7600 91.0500 2313.7600 93.0500 ;
        RECT 2552.2200 91.0500 2554.2200 93.0500 ;
        RECT 2792.6800 91.0500 2794.6800 93.0500 ;
        RECT 3033.1400 91.0500 3035.1400 93.0500 ;
        RECT 3273.6000 91.0500 3275.6000 93.0500 ;
        RECT 3514.0600 91.0500 3516.0600 93.0500 ;
        RECT 3754.5200 91.0500 3756.5200 93.0500 ;
        RECT 388.0800 3888.9100 390.0800 3890.9100 ;
        RECT 628.5400 3888.9100 630.5400 3890.9100 ;
        RECT 869.0000 3888.9100 871.0000 3890.9100 ;
        RECT 1109.4600 3888.9100 1111.4600 3890.9100 ;
        RECT 1349.9200 3888.9100 1351.9200 3890.9100 ;
        RECT 1590.3800 3888.9100 1592.3800 3890.9100 ;
        RECT 1830.8400 3888.9100 1832.8400 3890.9100 ;
        RECT 2071.3000 3888.9100 2073.3000 3890.9100 ;
        RECT 2311.7600 3888.9100 2313.7600 3890.9100 ;
        RECT 2552.2200 3888.9100 2554.2200 3890.9100 ;
        RECT 2792.6800 3888.9100 2794.6800 3890.9100 ;
        RECT 3033.1400 3888.9100 3035.1400 3890.9100 ;
        RECT 3273.6000 3888.9100 3275.6000 3890.9100 ;
        RECT 3514.0600 3888.9100 3516.0600 3890.9100 ;
        RECT 3754.5200 3888.9100 3756.5200 3890.9100 ;
      LAYER met5 ;
        RECT 157.0800 133.2400 3815.9800 135.2400 ;
        RECT 2.0000 82.9800 3766.0800 84.9800 ;
        RECT 2.0000 2.0000 3928.2400 6.0000 ;
        RECT 157.0800 383.0800 3815.9800 385.0800 ;
        RECT 157.0800 632.9200 3815.9800 634.9200 ;
        RECT 157.0800 882.7600 3815.9800 884.7600 ;
        RECT 157.0800 1882.1200 3815.9800 1884.1200 ;
        RECT 157.0800 1632.2800 3815.9800 1634.2800 ;
        RECT 157.0800 1382.4400 3815.9800 1384.4400 ;
        RECT 157.0800 1132.6000 3815.9800 1134.6000 ;
        RECT 2.0000 133.5000 159.0800 135.5000 ;
        RECT 389.0800 91.0500 399.6400 93.0500 ;
        RECT 2.0000 383.3400 159.0800 385.3400 ;
        RECT 121.1800 369.3400 159.0800 371.3400 ;
        RECT 629.5400 91.0500 640.1000 93.0500 ;
        RECT 870.0000 91.0500 880.5600 93.0500 ;
        RECT 121.1800 619.1800 159.0800 621.1800 ;
        RECT 2.0000 633.1800 159.0800 635.1800 ;
        RECT 121.1800 869.0200 159.0800 871.0200 ;
        RECT 2.0000 883.0200 159.0800 885.0200 ;
        RECT 1110.4600 91.0500 1121.0200 93.0500 ;
        RECT 1350.9200 91.0500 1361.4800 93.0500 ;
        RECT 1591.3800 91.0500 1601.9400 93.0500 ;
        RECT 1831.8400 91.0500 1842.4000 93.0500 ;
        RECT 121.1800 1118.8600 159.0800 1120.8600 ;
        RECT 2.0000 1132.8600 159.0800 1134.8600 ;
        RECT 121.1800 1368.7000 159.0800 1370.7000 ;
        RECT 2.0000 1382.7000 159.0800 1384.7000 ;
        RECT 121.1800 1618.5400 159.0800 1620.5400 ;
        RECT 2.0000 1632.5400 159.0800 1634.5400 ;
        RECT 121.1800 1868.3800 159.0800 1870.3800 ;
        RECT 2.0000 1882.3800 159.0800 1884.3800 ;
        RECT 2072.3000 91.0500 2082.8600 93.0500 ;
        RECT 2312.7600 91.0500 2323.3200 93.0500 ;
        RECT 2553.2200 91.0500 2563.7800 93.0500 ;
        RECT 2793.6800 91.0500 2804.2400 93.0500 ;
        RECT 3034.1400 91.0500 3044.7000 93.0500 ;
        RECT 3274.6000 91.0500 3285.1600 93.0500 ;
        RECT 3515.0600 91.0500 3525.6200 93.0500 ;
        RECT 3755.5200 91.0500 3766.0800 93.0500 ;
        RECT 2.0000 3924.0600 3928.2400 3928.0600 ;
        RECT 157.0800 2131.9600 3815.9800 2133.9600 ;
        RECT 157.0800 2381.8000 3815.9800 2383.8000 ;
        RECT 157.0800 2631.6400 3815.9800 2633.6400 ;
        RECT 157.0800 2881.4800 3815.9800 2883.4800 ;
        RECT 157.0800 3131.3200 3815.9800 3133.3200 ;
        RECT 157.0800 3381.1600 3815.9800 3383.1600 ;
        RECT 157.0800 3631.0000 3815.9800 3633.0000 ;
        RECT 157.0800 3880.8400 3766.0800 3882.8400 ;
        RECT 121.1800 2118.2200 159.0800 2120.2200 ;
        RECT 2.0000 2132.2200 159.0800 2134.2200 ;
        RECT 121.1800 2368.0600 159.0800 2370.0600 ;
        RECT 2.0000 2382.0600 159.0800 2384.0600 ;
        RECT 121.1800 2617.9000 159.0800 2619.9000 ;
        RECT 2.0000 2631.9000 159.0800 2633.9000 ;
        RECT 121.1800 2867.7400 159.0800 2869.7400 ;
        RECT 2.0000 2881.7400 159.0800 2883.7400 ;
        RECT 2.0000 3131.5800 159.0800 3133.5800 ;
        RECT 121.1800 3117.5800 159.0800 3119.5800 ;
        RECT 121.1800 3367.4200 159.0800 3369.4200 ;
        RECT 2.0000 3381.4200 159.0800 3383.4200 ;
        RECT 121.1800 3617.2600 159.0800 3619.2600 ;
        RECT 2.0000 3631.2600 159.0800 3633.2600 ;
        RECT 2.0000 3867.1000 159.0800 3869.1000 ;
        RECT 389.0800 3888.9100 399.6400 3890.9100 ;
        RECT 629.5400 3888.9100 640.1000 3890.9100 ;
        RECT 870.0000 3888.9100 880.5600 3890.9100 ;
        RECT 1110.4600 3888.9100 1121.0200 3890.9100 ;
        RECT 1350.9200 3888.9100 1361.4800 3890.9100 ;
        RECT 1591.3800 3888.9100 1601.9400 3890.9100 ;
        RECT 1831.8400 3888.9100 1842.4000 3890.9100 ;
        RECT 2072.3000 3888.9100 2082.8600 3890.9100 ;
        RECT 2312.7600 3888.9100 2323.3200 3890.9100 ;
        RECT 2553.2200 3888.9100 2563.7800 3890.9100 ;
        RECT 2793.6800 3888.9100 2804.2400 3890.9100 ;
        RECT 3034.1400 3888.9100 3044.7000 3890.9100 ;
        RECT 3274.6000 3888.9100 3285.1600 3890.9100 ;
        RECT 3515.0600 3888.9100 3525.6200 3890.9100 ;
        RECT 3755.5200 3888.9100 3766.0800 3890.9100 ;
        RECT 157.0800 133.2400 159.0800 135.5000 ;
        RECT 388.0800 91.0500 390.0800 93.0500 ;
        RECT 157.0800 383.0800 159.0800 385.3400 ;
        RECT 628.5400 91.0500 630.5400 93.0500 ;
        RECT 869.0000 91.0500 871.0000 93.0500 ;
        RECT 157.0800 632.9200 159.0800 635.1800 ;
        RECT 157.0800 882.7600 159.0800 885.0200 ;
        RECT 1109.4600 91.0500 1111.4600 93.0500 ;
        RECT 1349.9200 91.0500 1351.9200 93.0500 ;
        RECT 1590.3800 91.0500 1592.3800 93.0500 ;
        RECT 1830.8400 91.0500 1832.8400 93.0500 ;
        RECT 157.0800 1132.6000 159.0800 1134.8600 ;
        RECT 157.0800 1382.4400 159.0800 1384.7000 ;
        RECT 157.0800 1632.2800 159.0800 1634.5400 ;
        RECT 157.0800 1882.1200 159.0800 1884.3800 ;
        RECT 2071.3000 91.0500 2073.3000 93.0500 ;
        RECT 2311.7600 91.0500 2313.7600 93.0500 ;
        RECT 2552.2200 91.0500 2554.2200 93.0500 ;
        RECT 2792.6800 91.0500 2794.6800 93.0500 ;
        RECT 3033.1400 91.0500 3035.1400 93.0500 ;
        RECT 3273.6000 91.0500 3275.6000 93.0500 ;
        RECT 3514.0600 91.0500 3516.0600 93.0500 ;
        RECT 3754.5200 91.0500 3756.5200 93.0500 ;
        RECT 157.0800 2131.9600 159.0800 2134.2200 ;
        RECT 157.0800 2381.8000 159.0800 2384.0600 ;
        RECT 157.0800 2631.6400 159.0800 2633.9000 ;
        RECT 157.0800 2881.4800 159.0800 2883.7400 ;
        RECT 157.0800 3131.3200 159.0800 3133.5800 ;
        RECT 157.0800 3381.1600 159.0800 3383.4200 ;
        RECT 157.0800 3631.0000 159.0800 3633.2600 ;
        RECT 388.0800 3888.9100 390.0800 3890.9100 ;
        RECT 628.5400 3888.9100 630.5400 3890.9100 ;
        RECT 869.0000 3888.9100 871.0000 3890.9100 ;
        RECT 1109.4600 3888.9100 1111.4600 3890.9100 ;
        RECT 1349.9200 3888.9100 1351.9200 3890.9100 ;
        RECT 1590.3800 3888.9100 1592.3800 3890.9100 ;
        RECT 1830.8400 3888.9100 1832.8400 3890.9100 ;
        RECT 2071.3000 3888.9100 2073.3000 3890.9100 ;
        RECT 2311.7600 3888.9100 2313.7600 3890.9100 ;
        RECT 2552.2200 3888.9100 2554.2200 3890.9100 ;
        RECT 2792.6800 3888.9100 2794.6800 3890.9100 ;
        RECT 3033.1400 3888.9100 3035.1400 3890.9100 ;
        RECT 3273.6000 3888.9100 3275.6000 3890.9100 ;
        RECT 3514.0600 3888.9100 3516.0600 3890.9100 ;
        RECT 3754.5200 3888.9100 3756.5200 3890.9100 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 8.0000 8.0000 12.0000 3922.0600 ;
        RECT 117.1800 129.5000 119.1800 3629.2600 ;
        RECT 161.0800 129.5000 163.0800 3629.2600 ;
        RECT 401.6400 78.9800 403.6400 3922.0600 ;
        RECT 642.1000 78.9800 644.1000 3922.0600 ;
        RECT 882.5600 78.9800 884.5600 3922.0600 ;
        RECT 1844.4000 78.9800 1846.4000 3922.0600 ;
        RECT 1123.0200 78.9800 1125.0200 3922.0600 ;
        RECT 1363.4800 78.9800 1365.4800 3922.0600 ;
        RECT 1603.9400 78.9800 1605.9400 3922.0600 ;
        RECT 2806.2400 78.9800 2808.2400 3922.0600 ;
        RECT 2565.7800 78.9800 2567.7800 3922.0600 ;
        RECT 2325.3200 78.9800 2327.3200 3922.0600 ;
        RECT 2084.8600 78.9800 2086.8600 3922.0600 ;
        RECT 3778.0800 1878.1200 3780.0800 2117.9600 ;
        RECT 3817.9800 1878.1200 3819.9800 2117.9600 ;
        RECT 3768.0800 78.9800 3770.0800 3922.0600 ;
        RECT 3527.6200 78.9800 3529.6200 3922.0600 ;
        RECT 3287.1600 78.9800 3289.1600 3922.0600 ;
        RECT 3046.7000 78.9800 3048.7000 3922.0600 ;
        RECT 3918.2400 8.0000 3922.2400 3922.0600 ;
        RECT 161.1800 78.9800 163.1800 119.2400 ;
        RECT 161.1800 88.0500 168.7400 90.0500 ;
        RECT 161.0800 139.1700 168.2400 141.1700 ;
        RECT 152.0050 140.4300 154.6750 141.9300 ;
        RECT 161.0800 129.2400 163.0800 131.5000 ;
        RECT 401.6400 88.0500 409.2000 90.0500 ;
        RECT 401.6400 139.1700 408.7000 141.1700 ;
        RECT 161.0800 389.0100 168.2400 391.0100 ;
        RECT 152.0050 390.2700 154.6750 391.7700 ;
        RECT 401.6400 389.0100 408.7000 391.0100 ;
        RECT 642.1000 88.0500 649.6600 90.0500 ;
        RECT 642.1000 139.1700 649.1600 141.1700 ;
        RECT 882.5600 88.0500 890.1200 90.0500 ;
        RECT 882.5600 139.1700 889.6200 141.1700 ;
        RECT 642.1000 389.0100 649.1600 391.0100 ;
        RECT 882.5600 389.0100 889.6200 391.0100 ;
        RECT 161.0800 638.8500 168.2400 640.8500 ;
        RECT 152.0050 640.1100 154.6750 641.6100 ;
        RECT 401.6400 638.8500 408.7000 640.8500 ;
        RECT 161.0800 888.6900 168.2400 890.6900 ;
        RECT 152.0050 889.9500 154.6750 891.4500 ;
        RECT 401.6400 888.6900 408.7000 890.6900 ;
        RECT 642.1000 638.8500 649.1600 640.8500 ;
        RECT 882.5600 638.8500 889.6200 640.8500 ;
        RECT 642.1000 888.6900 649.1600 890.6900 ;
        RECT 882.5600 888.6900 889.6200 890.6900 ;
        RECT 1123.0200 88.0500 1130.5800 90.0500 ;
        RECT 1123.0200 139.1700 1130.0800 141.1700 ;
        RECT 1363.4800 88.0500 1371.0400 90.0500 ;
        RECT 1363.4800 139.1700 1370.5400 141.1700 ;
        RECT 1123.0200 389.0100 1130.0800 391.0100 ;
        RECT 1363.4800 389.0100 1370.5400 391.0100 ;
        RECT 1603.9400 88.0500 1611.5000 90.0500 ;
        RECT 1603.9400 139.1700 1611.0000 141.1700 ;
        RECT 1844.4000 88.0500 1851.9600 90.0500 ;
        RECT 1844.4000 139.1700 1851.4600 141.1700 ;
        RECT 1603.9400 389.0100 1611.0000 391.0100 ;
        RECT 1844.4000 389.0100 1851.4600 391.0100 ;
        RECT 1363.4800 638.8500 1370.5400 640.8500 ;
        RECT 1123.0200 638.8500 1130.0800 640.8500 ;
        RECT 1123.0200 888.6900 1130.0800 890.6900 ;
        RECT 1363.4800 888.6900 1370.5400 890.6900 ;
        RECT 1603.9400 638.8500 1611.0000 640.8500 ;
        RECT 1844.4000 638.8500 1851.4600 640.8500 ;
        RECT 1603.9400 888.6900 1611.0000 890.6900 ;
        RECT 1844.4000 888.6900 1851.4600 890.6900 ;
        RECT 161.0800 1138.5300 168.2400 1140.5300 ;
        RECT 152.0050 1139.7900 154.6750 1141.2900 ;
        RECT 401.6400 1138.5300 408.7000 1140.5300 ;
        RECT 161.0800 1388.3700 168.2400 1390.3700 ;
        RECT 152.0050 1389.6300 154.6750 1391.1300 ;
        RECT 401.6400 1388.3700 408.7000 1390.3700 ;
        RECT 642.1000 1138.5300 649.1600 1140.5300 ;
        RECT 882.5600 1138.5300 889.6200 1140.5300 ;
        RECT 642.1000 1388.3700 649.1600 1390.3700 ;
        RECT 882.5600 1388.3700 889.6200 1390.3700 ;
        RECT 161.0800 1638.2100 168.2400 1640.2100 ;
        RECT 152.0050 1639.4700 154.6750 1640.9700 ;
        RECT 401.6400 1638.2100 408.7000 1640.2100 ;
        RECT 161.0800 1888.0500 168.2400 1890.0500 ;
        RECT 152.0050 1889.3100 154.6750 1890.8100 ;
        RECT 401.6400 1888.0500 408.7000 1890.0500 ;
        RECT 642.1000 1638.2100 649.1600 1640.2100 ;
        RECT 882.5600 1638.2100 889.6200 1640.2100 ;
        RECT 882.5600 1888.0500 889.6200 1890.0500 ;
        RECT 642.1000 1888.0500 649.1600 1890.0500 ;
        RECT 1123.0200 1138.5300 1130.0800 1140.5300 ;
        RECT 1363.4800 1138.5300 1370.5400 1140.5300 ;
        RECT 1363.4800 1388.3700 1370.5400 1390.3700 ;
        RECT 1123.0200 1388.3700 1130.0800 1390.3700 ;
        RECT 1603.9400 1138.5300 1611.0000 1140.5300 ;
        RECT 1844.4000 1138.5300 1851.4600 1140.5300 ;
        RECT 1603.9400 1388.3700 1611.0000 1390.3700 ;
        RECT 1844.4000 1388.3700 1851.4600 1390.3700 ;
        RECT 1123.0200 1638.2100 1130.0800 1640.2100 ;
        RECT 1363.4800 1638.2100 1370.5400 1640.2100 ;
        RECT 1363.4800 1888.0500 1370.5400 1890.0500 ;
        RECT 1123.0200 1888.0500 1130.0800 1890.0500 ;
        RECT 1603.9400 1638.2100 1611.0000 1640.2100 ;
        RECT 1844.4000 1638.2100 1851.4600 1640.2100 ;
        RECT 1603.9400 1888.0500 1611.0000 1890.0500 ;
        RECT 1844.4000 1888.0500 1851.4600 1890.0500 ;
        RECT 3817.9800 878.7600 3819.9800 1118.6000 ;
        RECT 3778.0800 878.7600 3780.0800 1118.6000 ;
        RECT 2084.8600 88.0500 2092.4200 90.0500 ;
        RECT 2084.8600 139.1700 2091.9200 141.1700 ;
        RECT 2325.3200 88.0500 2332.8800 90.0500 ;
        RECT 2325.3200 139.1700 2332.3800 141.1700 ;
        RECT 2084.8600 389.0100 2091.9200 391.0100 ;
        RECT 2325.3200 389.0100 2332.3800 391.0100 ;
        RECT 2565.7800 88.0500 2573.3400 90.0500 ;
        RECT 2565.7800 139.1700 2572.8400 141.1700 ;
        RECT 2806.2400 88.0500 2813.8000 90.0500 ;
        RECT 2806.2400 139.1700 2813.3000 141.1700 ;
        RECT 2806.2400 389.0100 2813.3000 391.0100 ;
        RECT 2565.7800 389.0100 2572.8400 391.0100 ;
        RECT 2325.3200 638.8500 2332.3800 640.8500 ;
        RECT 2084.8600 638.8500 2091.9200 640.8500 ;
        RECT 2084.8600 888.6900 2091.9200 890.6900 ;
        RECT 2325.3200 888.6900 2332.3800 890.6900 ;
        RECT 2806.2400 638.8500 2813.3000 640.8500 ;
        RECT 2565.7800 638.8500 2572.8400 640.8500 ;
        RECT 2806.2400 888.6900 2813.3000 890.6900 ;
        RECT 2565.7800 888.6900 2572.8400 890.6900 ;
        RECT 3817.9800 379.0800 3819.9800 618.9200 ;
        RECT 3778.0800 379.0800 3780.0800 618.9200 ;
        RECT 3046.7000 88.0500 3054.2600 90.0500 ;
        RECT 3046.7000 139.1700 3053.7600 141.1700 ;
        RECT 3287.1600 88.0500 3294.7200 90.0500 ;
        RECT 3287.1600 139.1700 3294.2200 141.1700 ;
        RECT 3046.7000 389.0100 3053.7600 391.0100 ;
        RECT 3287.1600 389.0100 3294.2200 391.0100 ;
        RECT 3817.9800 129.2400 3819.9800 369.0800 ;
        RECT 3778.0800 129.2400 3780.0800 369.0800 ;
        RECT 3527.6200 139.1700 3534.6800 141.1700 ;
        RECT 3527.6200 88.0500 3535.1800 90.0500 ;
        RECT 3778.0800 140.1700 3783.8200 141.6700 ;
        RECT 3527.6200 389.0100 3534.6800 391.0100 ;
        RECT 3778.0800 390.0100 3783.8200 391.5100 ;
        RECT 3046.7000 638.8500 3053.7600 640.8500 ;
        RECT 3287.1600 638.8500 3294.2200 640.8500 ;
        RECT 3046.7000 888.6900 3053.7600 890.6900 ;
        RECT 3287.1600 888.6900 3294.2200 890.6900 ;
        RECT 3778.0800 628.9200 3780.0800 868.7600 ;
        RECT 3817.9800 628.9200 3819.9800 868.7600 ;
        RECT 3527.6200 638.8500 3534.6800 640.8500 ;
        RECT 3778.0800 639.8500 3783.8200 641.3500 ;
        RECT 3527.6200 888.6900 3534.6800 890.6900 ;
        RECT 3778.0800 889.6900 3783.8200 891.1900 ;
        RECT 2084.8600 1138.5300 2091.9200 1140.5300 ;
        RECT 2325.3200 1138.5300 2332.3800 1140.5300 ;
        RECT 2325.3200 1388.3700 2332.3800 1390.3700 ;
        RECT 2084.8600 1388.3700 2091.9200 1390.3700 ;
        RECT 2806.2400 1138.5300 2813.3000 1140.5300 ;
        RECT 2565.7800 1138.5300 2572.8400 1140.5300 ;
        RECT 2806.2400 1388.3700 2813.3000 1390.3700 ;
        RECT 2565.7800 1388.3700 2572.8400 1390.3700 ;
        RECT 2084.8600 1638.2100 2091.9200 1640.2100 ;
        RECT 2325.3200 1638.2100 2332.3800 1640.2100 ;
        RECT 2325.3200 1888.0500 2332.3800 1890.0500 ;
        RECT 2084.8600 1888.0500 2091.9200 1890.0500 ;
        RECT 2806.2400 1638.2100 2813.3000 1640.2100 ;
        RECT 2565.7800 1638.2100 2572.8400 1640.2100 ;
        RECT 2806.2400 1888.0500 2813.3000 1890.0500 ;
        RECT 2565.7800 1888.0500 2572.8400 1890.0500 ;
        RECT 3817.9800 1378.4400 3819.9800 1618.2800 ;
        RECT 3778.0800 1378.4400 3780.0800 1618.2800 ;
        RECT 3046.7000 1138.5300 3053.7600 1140.5300 ;
        RECT 3287.1600 1138.5300 3294.2200 1140.5300 ;
        RECT 3287.1600 1388.3700 3294.2200 1390.3700 ;
        RECT 3046.7000 1388.3700 3053.7600 1390.3700 ;
        RECT 3778.0800 1128.6000 3780.0800 1368.4400 ;
        RECT 3817.9800 1128.6000 3819.9800 1368.4400 ;
        RECT 3527.6200 1138.5300 3534.6800 1140.5300 ;
        RECT 3778.0800 1139.5300 3783.8200 1141.0300 ;
        RECT 3527.6200 1388.3700 3534.6800 1390.3700 ;
        RECT 3778.0800 1389.3700 3783.8200 1390.8700 ;
        RECT 3287.1600 1638.2100 3294.2200 1640.2100 ;
        RECT 3046.7000 1638.2100 3053.7600 1640.2100 ;
        RECT 3287.1600 1888.0500 3294.2200 1890.0500 ;
        RECT 3046.7000 1888.0500 3053.7600 1890.0500 ;
        RECT 3778.0800 1628.2800 3780.0800 1868.1200 ;
        RECT 3817.9800 1628.2800 3819.9800 1868.1200 ;
        RECT 3527.6200 1638.2100 3534.6800 1640.2100 ;
        RECT 3778.0800 1639.2100 3783.8200 1640.7100 ;
        RECT 3527.6200 1888.0500 3534.6800 1890.0500 ;
        RECT 3778.0800 1889.0500 3783.8200 1890.5500 ;
        RECT 161.0800 2137.8900 168.2400 2139.8900 ;
        RECT 152.0050 2139.1500 154.6750 2140.6500 ;
        RECT 401.6400 2137.8900 408.7000 2139.8900 ;
        RECT 161.0800 2387.7300 168.2400 2389.7300 ;
        RECT 152.0050 2388.9900 154.6750 2390.4900 ;
        RECT 401.6400 2387.7300 408.7000 2389.7300 ;
        RECT 882.5600 2137.8900 889.6200 2139.8900 ;
        RECT 642.1000 2137.8900 649.1600 2139.8900 ;
        RECT 882.5600 2387.7300 889.6200 2389.7300 ;
        RECT 642.1000 2387.7300 649.1600 2389.7300 ;
        RECT 161.0800 2637.5700 168.2400 2639.5700 ;
        RECT 152.0050 2638.8300 154.6750 2640.3300 ;
        RECT 401.6400 2637.5700 408.7000 2639.5700 ;
        RECT 161.0800 2887.4100 168.2400 2889.4100 ;
        RECT 152.0050 2888.6700 154.6750 2890.1700 ;
        RECT 401.6400 2887.4100 408.7000 2889.4100 ;
        RECT 882.5600 2637.5700 889.6200 2639.5700 ;
        RECT 642.1000 2637.5700 649.1600 2639.5700 ;
        RECT 882.5600 2887.4100 889.6200 2889.4100 ;
        RECT 642.1000 2887.4100 649.1600 2889.4100 ;
        RECT 1363.4800 2137.8900 1370.5400 2139.8900 ;
        RECT 1123.0200 2137.8900 1130.0800 2139.8900 ;
        RECT 1123.0200 2387.7300 1130.0800 2389.7300 ;
        RECT 1363.4800 2387.7300 1370.5400 2389.7300 ;
        RECT 1603.9400 2137.8900 1611.0000 2139.8900 ;
        RECT 1844.4000 2137.8900 1851.4600 2139.8900 ;
        RECT 1603.9400 2387.7300 1611.0000 2389.7300 ;
        RECT 1844.4000 2387.7300 1851.4600 2389.7300 ;
        RECT 1363.4800 2637.5700 1370.5400 2639.5700 ;
        RECT 1123.0200 2637.5700 1130.0800 2639.5700 ;
        RECT 1123.0200 2887.4100 1130.0800 2889.4100 ;
        RECT 1363.4800 2887.4100 1370.5400 2889.4100 ;
        RECT 1603.9400 2637.5700 1611.0000 2639.5700 ;
        RECT 1844.4000 2637.5700 1851.4600 2639.5700 ;
        RECT 1603.9400 2887.4100 1611.0000 2889.4100 ;
        RECT 1844.4000 2887.4100 1851.4600 2889.4100 ;
        RECT 161.0800 3137.2500 168.2400 3139.2500 ;
        RECT 152.0050 3138.5100 154.6750 3140.0100 ;
        RECT 401.6400 3137.2500 408.7000 3139.2500 ;
        RECT 161.0800 3387.0900 168.2400 3389.0900 ;
        RECT 152.0050 3388.3500 154.6750 3389.8500 ;
        RECT 401.6400 3387.0900 408.7000 3389.0900 ;
        RECT 642.1000 3137.2500 649.1600 3139.2500 ;
        RECT 882.5600 3137.2500 889.6200 3139.2500 ;
        RECT 642.1000 3387.0900 649.1600 3389.0900 ;
        RECT 882.5600 3387.0900 889.6200 3389.0900 ;
        RECT 117.1800 3627.2600 119.1800 3922.0600 ;
        RECT 161.0800 3627.2600 163.0800 3922.0600 ;
        RECT 161.0800 3636.9300 168.2400 3638.9300 ;
        RECT 152.0050 3638.1900 154.6750 3639.6900 ;
        RECT 401.6400 3636.9300 408.7000 3638.9300 ;
        RECT 161.0800 3910.8400 168.7400 3912.8400 ;
        RECT 401.6400 3910.8400 409.2000 3912.8400 ;
        RECT 401.6400 3882.8400 403.6400 3922.0600 ;
        RECT 642.1000 3636.9300 649.1600 3638.9300 ;
        RECT 882.5600 3636.9300 889.6200 3638.9300 ;
        RECT 642.1000 3882.8400 644.1000 3922.0600 ;
        RECT 642.1000 3910.8400 649.6600 3912.8400 ;
        RECT 882.5600 3882.8400 884.5600 3922.0600 ;
        RECT 882.5600 3910.8400 890.1200 3912.8400 ;
        RECT 1123.0200 3137.2500 1130.0800 3139.2500 ;
        RECT 1363.4800 3137.2500 1370.5400 3139.2500 ;
        RECT 1123.0200 3387.0900 1130.0800 3389.0900 ;
        RECT 1363.4800 3387.0900 1370.5400 3389.0900 ;
        RECT 1603.9400 3137.2500 1611.0000 3139.2500 ;
        RECT 1844.4000 3137.2500 1851.4600 3139.2500 ;
        RECT 1603.9400 3387.0900 1611.0000 3389.0900 ;
        RECT 1844.4000 3387.0900 1851.4600 3389.0900 ;
        RECT 1123.0200 3636.9300 1130.0800 3638.9300 ;
        RECT 1363.4800 3636.9300 1370.5400 3638.9300 ;
        RECT 1123.0200 3882.8400 1125.0200 3922.0600 ;
        RECT 1123.0200 3910.8400 1130.5800 3912.8400 ;
        RECT 1363.4800 3882.8400 1365.4800 3922.0600 ;
        RECT 1363.4800 3910.8400 1371.0400 3912.8400 ;
        RECT 1844.4000 3636.9300 1851.4600 3638.9300 ;
        RECT 1603.9400 3636.9300 1611.0000 3638.9300 ;
        RECT 1603.9400 3882.8400 1605.9400 3922.0600 ;
        RECT 1603.9400 3910.8400 1611.5000 3912.8400 ;
        RECT 1844.4000 3882.8400 1846.4000 3922.0600 ;
        RECT 1844.4000 3910.8400 1851.9600 3912.8400 ;
        RECT 3817.9800 2877.4800 3819.9800 3117.3200 ;
        RECT 3778.0800 2877.4800 3780.0800 3117.3200 ;
        RECT 2084.8600 2137.8900 2091.9200 2139.8900 ;
        RECT 2325.3200 2137.8900 2332.3800 2139.8900 ;
        RECT 2325.3200 2387.7300 2332.3800 2389.7300 ;
        RECT 2084.8600 2387.7300 2091.9200 2389.7300 ;
        RECT 2806.2400 2137.8900 2813.3000 2139.8900 ;
        RECT 2565.7800 2137.8900 2572.8400 2139.8900 ;
        RECT 2806.2400 2387.7300 2813.3000 2389.7300 ;
        RECT 2565.7800 2387.7300 2572.8400 2389.7300 ;
        RECT 2325.3200 2637.5700 2332.3800 2639.5700 ;
        RECT 2084.8600 2637.5700 2091.9200 2639.5700 ;
        RECT 2084.8600 2887.4100 2091.9200 2889.4100 ;
        RECT 2325.3200 2887.4100 2332.3800 2889.4100 ;
        RECT 2806.2400 2637.5700 2813.3000 2639.5700 ;
        RECT 2565.7800 2637.5700 2572.8400 2639.5700 ;
        RECT 2806.2400 2887.4100 2813.3000 2889.4100 ;
        RECT 2565.7800 2887.4100 2572.8400 2889.4100 ;
        RECT 3817.9800 2377.8000 3819.9800 2617.6400 ;
        RECT 3778.0800 2377.8000 3780.0800 2617.6400 ;
        RECT 3287.1600 2137.8900 3294.2200 2139.8900 ;
        RECT 3046.7000 2137.8900 3053.7600 2139.8900 ;
        RECT 3287.1600 2387.7300 3294.2200 2389.7300 ;
        RECT 3046.7000 2387.7300 3053.7600 2389.7300 ;
        RECT 3778.0800 2127.9600 3780.0800 2367.8000 ;
        RECT 3817.9800 2127.9600 3819.9800 2367.8000 ;
        RECT 3527.6200 2137.8900 3534.6800 2139.8900 ;
        RECT 3778.0800 2138.8900 3783.8200 2140.3900 ;
        RECT 3527.6200 2387.7300 3534.6800 2389.7300 ;
        RECT 3778.0800 2388.7300 3783.8200 2390.2300 ;
        RECT 3287.1600 2637.5700 3294.2200 2639.5700 ;
        RECT 3046.7000 2637.5700 3053.7600 2639.5700 ;
        RECT 3287.1600 2887.4100 3294.2200 2889.4100 ;
        RECT 3046.7000 2887.4100 3053.7600 2889.4100 ;
        RECT 3778.0800 2627.6400 3780.0800 2867.4800 ;
        RECT 3817.9800 2627.6400 3819.9800 2867.4800 ;
        RECT 3527.6200 2637.5700 3534.6800 2639.5700 ;
        RECT 3778.0800 2638.5700 3783.8200 2640.0700 ;
        RECT 3527.6200 2887.4100 3534.6800 2889.4100 ;
        RECT 3778.0800 2888.4100 3783.8200 2889.9100 ;
        RECT 2325.3200 3137.2500 2332.3800 3139.2500 ;
        RECT 2084.8600 3137.2500 2091.9200 3139.2500 ;
        RECT 2084.8600 3387.0900 2091.9200 3389.0900 ;
        RECT 2325.3200 3387.0900 2332.3800 3389.0900 ;
        RECT 2806.2400 3137.2500 2813.3000 3139.2500 ;
        RECT 2565.7800 3137.2500 2572.8400 3139.2500 ;
        RECT 2806.2400 3387.0900 2813.3000 3389.0900 ;
        RECT 2565.7800 3387.0900 2572.8400 3389.0900 ;
        RECT 2084.8600 3636.9300 2091.9200 3638.9300 ;
        RECT 2325.3200 3636.9300 2332.3800 3638.9300 ;
        RECT 2084.8600 3882.8400 2086.8600 3922.0600 ;
        RECT 2084.8600 3910.8400 2092.4200 3912.8400 ;
        RECT 2325.3200 3882.8400 2327.3200 3922.0600 ;
        RECT 2325.3200 3910.8400 2332.8800 3912.8400 ;
        RECT 2806.2400 3636.9300 2813.3000 3638.9300 ;
        RECT 2565.7800 3882.8400 2567.7800 3922.0600 ;
        RECT 2565.7800 3910.8400 2573.3400 3912.8400 ;
        RECT 2806.2400 3882.8400 2808.2400 3922.0600 ;
        RECT 2806.2400 3910.8400 2813.8000 3912.8400 ;
        RECT 3817.9800 3377.1600 3819.9800 3617.0000 ;
        RECT 3778.0800 3377.1600 3780.0800 3617.0000 ;
        RECT 3287.1600 3137.2500 3294.2200 3139.2500 ;
        RECT 3046.7000 3137.2500 3053.7600 3139.2500 ;
        RECT 3287.1600 3387.0900 3294.2200 3389.0900 ;
        RECT 3046.7000 3387.0900 3053.7600 3389.0900 ;
        RECT 3778.0800 3127.3200 3780.0800 3367.1600 ;
        RECT 3817.9800 3127.3200 3819.9800 3367.1600 ;
        RECT 3527.6200 3137.2500 3534.6800 3139.2500 ;
        RECT 3778.0800 3138.2500 3783.8200 3139.7500 ;
        RECT 3527.6200 3387.0900 3534.6800 3389.0900 ;
        RECT 3778.0800 3388.0900 3783.8200 3389.5900 ;
        RECT 3287.1600 3636.9300 3294.2200 3638.9300 ;
        RECT 3046.7000 3636.9300 3053.7600 3638.9300 ;
        RECT 3046.7000 3882.8400 3048.7000 3922.0600 ;
        RECT 3046.7000 3910.8400 3054.2600 3912.8400 ;
        RECT 3287.1600 3882.8400 3289.1600 3922.0600 ;
        RECT 3287.1600 3910.8400 3294.7200 3912.8400 ;
        RECT 3817.9800 3627.0000 3819.9800 3866.8400 ;
        RECT 3778.0800 3627.0000 3780.0800 3866.8400 ;
        RECT 3527.6200 3636.9300 3534.6800 3638.9300 ;
        RECT 3778.0800 3637.9300 3783.8200 3639.4300 ;
        RECT 3527.6200 3882.8400 3529.6200 3922.0600 ;
        RECT 3527.6200 3910.8400 3535.1800 3912.8400 ;
        RECT 3768.0800 3882.8400 3770.0800 3922.0600 ;
        RECT 167.7400 88.0500 169.7400 90.0500 ;
        RECT 166.7400 139.1700 169.7400 141.1700 ;
        RECT 408.2000 88.0500 410.2000 90.0500 ;
        RECT 407.2000 139.1700 410.2000 141.1700 ;
        RECT 166.7400 389.0100 169.7400 391.0100 ;
        RECT 407.2000 389.0100 410.2000 391.0100 ;
        RECT 648.6600 88.0500 650.6600 90.0500 ;
        RECT 647.6600 139.1700 650.6600 141.1700 ;
        RECT 889.1200 88.0500 891.1200 90.0500 ;
        RECT 888.1200 139.1700 891.1200 141.1700 ;
        RECT 647.6600 389.0100 650.6600 391.0100 ;
        RECT 888.1200 389.0100 891.1200 391.0100 ;
        RECT 166.7400 638.8500 169.7400 640.8500 ;
        RECT 407.2000 638.8500 410.2000 640.8500 ;
        RECT 166.7400 888.6900 169.7400 890.6900 ;
        RECT 407.2000 888.6900 410.2000 890.6900 ;
        RECT 647.6600 638.8500 650.6600 640.8500 ;
        RECT 888.1200 638.8500 891.1200 640.8500 ;
        RECT 647.6600 888.6900 650.6600 890.6900 ;
        RECT 888.1200 888.6900 891.1200 890.6900 ;
        RECT 1129.5800 88.0500 1131.5800 90.0500 ;
        RECT 1128.5800 139.1700 1131.5800 141.1700 ;
        RECT 1370.0400 88.0500 1372.0400 90.0500 ;
        RECT 1369.0400 139.1700 1372.0400 141.1700 ;
        RECT 1128.5800 389.0100 1131.5800 391.0100 ;
        RECT 1369.0400 389.0100 1372.0400 391.0100 ;
        RECT 1610.5000 88.0500 1612.5000 90.0500 ;
        RECT 1609.5000 139.1700 1612.5000 141.1700 ;
        RECT 1850.9600 88.0500 1852.9600 90.0500 ;
        RECT 1849.9600 139.1700 1852.9600 141.1700 ;
        RECT 1609.5000 389.0100 1612.5000 391.0100 ;
        RECT 1849.9600 389.0100 1852.9600 391.0100 ;
        RECT 1128.5800 638.8500 1131.5800 640.8500 ;
        RECT 1369.0400 638.8500 1372.0400 640.8500 ;
        RECT 1128.5800 888.6900 1131.5800 890.6900 ;
        RECT 1369.0400 888.6900 1372.0400 890.6900 ;
        RECT 1609.5000 638.8500 1612.5000 640.8500 ;
        RECT 1849.9600 638.8500 1852.9600 640.8500 ;
        RECT 1609.5000 888.6900 1612.5000 890.6900 ;
        RECT 1849.9600 888.6900 1852.9600 890.6900 ;
        RECT 166.7400 1138.5300 169.7400 1140.5300 ;
        RECT 407.2000 1138.5300 410.2000 1140.5300 ;
        RECT 166.7400 1388.3700 169.7400 1390.3700 ;
        RECT 407.2000 1388.3700 410.2000 1390.3700 ;
        RECT 647.6600 1138.5300 650.6600 1140.5300 ;
        RECT 888.1200 1138.5300 891.1200 1140.5300 ;
        RECT 647.6600 1388.3700 650.6600 1390.3700 ;
        RECT 888.1200 1388.3700 891.1200 1390.3700 ;
        RECT 166.7400 1638.2100 169.7400 1640.2100 ;
        RECT 407.2000 1638.2100 410.2000 1640.2100 ;
        RECT 166.7400 1888.0500 169.7400 1890.0500 ;
        RECT 407.2000 1888.0500 410.2000 1890.0500 ;
        RECT 647.6600 1638.2100 650.6600 1640.2100 ;
        RECT 888.1200 1638.2100 891.1200 1640.2100 ;
        RECT 647.6600 1888.0500 650.6600 1890.0500 ;
        RECT 888.1200 1888.0500 891.1200 1890.0500 ;
        RECT 1128.5800 1138.5300 1131.5800 1140.5300 ;
        RECT 1369.0400 1138.5300 1372.0400 1140.5300 ;
        RECT 1128.5800 1388.3700 1131.5800 1390.3700 ;
        RECT 1369.0400 1388.3700 1372.0400 1390.3700 ;
        RECT 1609.5000 1138.5300 1612.5000 1140.5300 ;
        RECT 1849.9600 1138.5300 1852.9600 1140.5300 ;
        RECT 1609.5000 1388.3700 1612.5000 1390.3700 ;
        RECT 1849.9600 1388.3700 1852.9600 1390.3700 ;
        RECT 1128.5800 1638.2100 1131.5800 1640.2100 ;
        RECT 1369.0400 1638.2100 1372.0400 1640.2100 ;
        RECT 1128.5800 1888.0500 1131.5800 1890.0500 ;
        RECT 1369.0400 1888.0500 1372.0400 1890.0500 ;
        RECT 1609.5000 1638.2100 1612.5000 1640.2100 ;
        RECT 1849.9600 1638.2100 1852.9600 1640.2100 ;
        RECT 1609.5000 1888.0500 1612.5000 1890.0500 ;
        RECT 1849.9600 1888.0500 1852.9600 1890.0500 ;
        RECT 2091.4200 88.0500 2093.4200 90.0500 ;
        RECT 2090.4200 139.1700 2093.4200 141.1700 ;
        RECT 2331.8800 88.0500 2333.8800 90.0500 ;
        RECT 2330.8800 139.1700 2333.8800 141.1700 ;
        RECT 2090.4200 389.0100 2093.4200 391.0100 ;
        RECT 2330.8800 389.0100 2333.8800 391.0100 ;
        RECT 2572.3400 88.0500 2574.3400 90.0500 ;
        RECT 2571.3400 139.1700 2574.3400 141.1700 ;
        RECT 2812.8000 88.0500 2814.8000 90.0500 ;
        RECT 2811.8000 139.1700 2814.8000 141.1700 ;
        RECT 2571.3400 389.0100 2574.3400 391.0100 ;
        RECT 2811.8000 389.0100 2814.8000 391.0100 ;
        RECT 2090.4200 638.8500 2093.4200 640.8500 ;
        RECT 2330.8800 638.8500 2333.8800 640.8500 ;
        RECT 2090.4200 888.6900 2093.4200 890.6900 ;
        RECT 2330.8800 888.6900 2333.8800 890.6900 ;
        RECT 2571.3400 638.8500 2574.3400 640.8500 ;
        RECT 2811.8000 638.8500 2814.8000 640.8500 ;
        RECT 2571.3400 888.6900 2574.3400 890.6900 ;
        RECT 2811.8000 888.6900 2814.8000 890.6900 ;
        RECT 3053.2600 88.0500 3055.2600 90.0500 ;
        RECT 3052.2600 139.1700 3055.2600 141.1700 ;
        RECT 3293.7200 88.0500 3295.7200 90.0500 ;
        RECT 3292.7200 139.1700 3295.7200 141.1700 ;
        RECT 3052.2600 389.0100 3055.2600 391.0100 ;
        RECT 3292.7200 389.0100 3295.7200 391.0100 ;
        RECT 3534.1800 88.0500 3536.1800 90.0500 ;
        RECT 3533.1800 139.1700 3536.1800 141.1700 ;
        RECT 3783.0700 140.1700 3784.5700 141.6700 ;
        RECT 3533.1800 389.0100 3536.1800 391.0100 ;
        RECT 3783.0700 390.0100 3784.5700 391.5100 ;
        RECT 3052.2600 638.8500 3055.2600 640.8500 ;
        RECT 3292.7200 638.8500 3295.7200 640.8500 ;
        RECT 3052.2600 888.6900 3055.2600 890.6900 ;
        RECT 3292.7200 888.6900 3295.7200 890.6900 ;
        RECT 3533.1800 638.8500 3536.1800 640.8500 ;
        RECT 3783.0700 639.8500 3784.5700 641.3500 ;
        RECT 3533.1800 888.6900 3536.1800 890.6900 ;
        RECT 3783.0700 889.6900 3784.5700 891.1900 ;
        RECT 2090.4200 1138.5300 2093.4200 1140.5300 ;
        RECT 2330.8800 1138.5300 2333.8800 1140.5300 ;
        RECT 2090.4200 1388.3700 2093.4200 1390.3700 ;
        RECT 2330.8800 1388.3700 2333.8800 1390.3700 ;
        RECT 2571.3400 1138.5300 2574.3400 1140.5300 ;
        RECT 2811.8000 1138.5300 2814.8000 1140.5300 ;
        RECT 2571.3400 1388.3700 2574.3400 1390.3700 ;
        RECT 2811.8000 1388.3700 2814.8000 1390.3700 ;
        RECT 2090.4200 1638.2100 2093.4200 1640.2100 ;
        RECT 2330.8800 1638.2100 2333.8800 1640.2100 ;
        RECT 2090.4200 1888.0500 2093.4200 1890.0500 ;
        RECT 2330.8800 1888.0500 2333.8800 1890.0500 ;
        RECT 2571.3400 1638.2100 2574.3400 1640.2100 ;
        RECT 2811.8000 1638.2100 2814.8000 1640.2100 ;
        RECT 2571.3400 1888.0500 2574.3400 1890.0500 ;
        RECT 2811.8000 1888.0500 2814.8000 1890.0500 ;
        RECT 3052.2600 1138.5300 3055.2600 1140.5300 ;
        RECT 3292.7200 1138.5300 3295.7200 1140.5300 ;
        RECT 3052.2600 1388.3700 3055.2600 1390.3700 ;
        RECT 3292.7200 1388.3700 3295.7200 1390.3700 ;
        RECT 3533.1800 1138.5300 3536.1800 1140.5300 ;
        RECT 3783.0700 1139.5300 3784.5700 1141.0300 ;
        RECT 3533.1800 1388.3700 3536.1800 1390.3700 ;
        RECT 3783.0700 1389.3700 3784.5700 1390.8700 ;
        RECT 3052.2600 1638.2100 3055.2600 1640.2100 ;
        RECT 3292.7200 1638.2100 3295.7200 1640.2100 ;
        RECT 3052.2600 1888.0500 3055.2600 1890.0500 ;
        RECT 3292.7200 1888.0500 3295.7200 1890.0500 ;
        RECT 3533.1800 1638.2100 3536.1800 1640.2100 ;
        RECT 3783.0700 1639.2100 3784.5700 1640.7100 ;
        RECT 3533.1800 1888.0500 3536.1800 1890.0500 ;
        RECT 3783.0700 1889.0500 3784.5700 1890.5500 ;
        RECT 166.7400 2137.8900 169.7400 2139.8900 ;
        RECT 407.2000 2137.8900 410.2000 2139.8900 ;
        RECT 166.7400 2387.7300 169.7400 2389.7300 ;
        RECT 407.2000 2387.7300 410.2000 2389.7300 ;
        RECT 647.6600 2137.8900 650.6600 2139.8900 ;
        RECT 888.1200 2137.8900 891.1200 2139.8900 ;
        RECT 647.6600 2387.7300 650.6600 2389.7300 ;
        RECT 888.1200 2387.7300 891.1200 2389.7300 ;
        RECT 166.7400 2637.5700 169.7400 2639.5700 ;
        RECT 407.2000 2637.5700 410.2000 2639.5700 ;
        RECT 166.7400 2887.4100 169.7400 2889.4100 ;
        RECT 407.2000 2887.4100 410.2000 2889.4100 ;
        RECT 647.6600 2637.5700 650.6600 2639.5700 ;
        RECT 888.1200 2637.5700 891.1200 2639.5700 ;
        RECT 647.6600 2887.4100 650.6600 2889.4100 ;
        RECT 888.1200 2887.4100 891.1200 2889.4100 ;
        RECT 1128.5800 2137.8900 1131.5800 2139.8900 ;
        RECT 1369.0400 2137.8900 1372.0400 2139.8900 ;
        RECT 1128.5800 2387.7300 1131.5800 2389.7300 ;
        RECT 1369.0400 2387.7300 1372.0400 2389.7300 ;
        RECT 1609.5000 2137.8900 1612.5000 2139.8900 ;
        RECT 1849.9600 2137.8900 1852.9600 2139.8900 ;
        RECT 1609.5000 2387.7300 1612.5000 2389.7300 ;
        RECT 1849.9600 2387.7300 1852.9600 2389.7300 ;
        RECT 1128.5800 2637.5700 1131.5800 2639.5700 ;
        RECT 1369.0400 2637.5700 1372.0400 2639.5700 ;
        RECT 1128.5800 2887.4100 1131.5800 2889.4100 ;
        RECT 1369.0400 2887.4100 1372.0400 2889.4100 ;
        RECT 1609.5000 2637.5700 1612.5000 2639.5700 ;
        RECT 1849.9600 2637.5700 1852.9600 2639.5700 ;
        RECT 1609.5000 2887.4100 1612.5000 2889.4100 ;
        RECT 1849.9600 2887.4100 1852.9600 2889.4100 ;
        RECT 166.7400 3137.2500 169.7400 3139.2500 ;
        RECT 407.2000 3137.2500 410.2000 3139.2500 ;
        RECT 166.7400 3387.0900 169.7400 3389.0900 ;
        RECT 407.2000 3387.0900 410.2000 3389.0900 ;
        RECT 647.6600 3137.2500 650.6600 3139.2500 ;
        RECT 888.1200 3137.2500 891.1200 3139.2500 ;
        RECT 647.6600 3387.0900 650.6600 3389.0900 ;
        RECT 888.1200 3387.0900 891.1200 3389.0900 ;
        RECT 166.7400 3636.9300 169.7400 3638.9300 ;
        RECT 407.2000 3636.9300 410.2000 3638.9300 ;
        RECT 167.7400 3910.8400 169.7400 3912.8400 ;
        RECT 408.2000 3910.8400 410.2000 3912.8400 ;
        RECT 647.6600 3636.9300 650.6600 3638.9300 ;
        RECT 888.1200 3636.9300 891.1200 3638.9300 ;
        RECT 648.6600 3910.8400 650.6600 3912.8400 ;
        RECT 889.1200 3910.8400 891.1200 3912.8400 ;
        RECT 1128.5800 3137.2500 1131.5800 3139.2500 ;
        RECT 1369.0400 3137.2500 1372.0400 3139.2500 ;
        RECT 1128.5800 3387.0900 1131.5800 3389.0900 ;
        RECT 1369.0400 3387.0900 1372.0400 3389.0900 ;
        RECT 1609.5000 3137.2500 1612.5000 3139.2500 ;
        RECT 1849.9600 3137.2500 1852.9600 3139.2500 ;
        RECT 1609.5000 3387.0900 1612.5000 3389.0900 ;
        RECT 1849.9600 3387.0900 1852.9600 3389.0900 ;
        RECT 1128.5800 3636.9300 1131.5800 3638.9300 ;
        RECT 1369.0400 3636.9300 1372.0400 3638.9300 ;
        RECT 1129.5800 3910.8400 1131.5800 3912.8400 ;
        RECT 1370.0400 3910.8400 1372.0400 3912.8400 ;
        RECT 1609.5000 3636.9300 1612.5000 3638.9300 ;
        RECT 1849.9600 3636.9300 1852.9600 3638.9300 ;
        RECT 1610.5000 3910.8400 1612.5000 3912.8400 ;
        RECT 1850.9600 3910.8400 1852.9600 3912.8400 ;
        RECT 2090.4200 2137.8900 2093.4200 2139.8900 ;
        RECT 2330.8800 2137.8900 2333.8800 2139.8900 ;
        RECT 2090.4200 2387.7300 2093.4200 2389.7300 ;
        RECT 2330.8800 2387.7300 2333.8800 2389.7300 ;
        RECT 2571.3400 2137.8900 2574.3400 2139.8900 ;
        RECT 2811.8000 2137.8900 2814.8000 2139.8900 ;
        RECT 2571.3400 2387.7300 2574.3400 2389.7300 ;
        RECT 2811.8000 2387.7300 2814.8000 2389.7300 ;
        RECT 2090.4200 2637.5700 2093.4200 2639.5700 ;
        RECT 2330.8800 2637.5700 2333.8800 2639.5700 ;
        RECT 2090.4200 2887.4100 2093.4200 2889.4100 ;
        RECT 2330.8800 2887.4100 2333.8800 2889.4100 ;
        RECT 2571.3400 2637.5700 2574.3400 2639.5700 ;
        RECT 2811.8000 2637.5700 2814.8000 2639.5700 ;
        RECT 2571.3400 2887.4100 2574.3400 2889.4100 ;
        RECT 2811.8000 2887.4100 2814.8000 2889.4100 ;
        RECT 3052.2600 2137.8900 3055.2600 2139.8900 ;
        RECT 3292.7200 2137.8900 3295.7200 2139.8900 ;
        RECT 3052.2600 2387.7300 3055.2600 2389.7300 ;
        RECT 3292.7200 2387.7300 3295.7200 2389.7300 ;
        RECT 3533.1800 2137.8900 3536.1800 2139.8900 ;
        RECT 3783.0700 2138.8900 3784.5700 2140.3900 ;
        RECT 3533.1800 2387.7300 3536.1800 2389.7300 ;
        RECT 3783.0700 2388.7300 3784.5700 2390.2300 ;
        RECT 3052.2600 2637.5700 3055.2600 2639.5700 ;
        RECT 3292.7200 2637.5700 3295.7200 2639.5700 ;
        RECT 3052.2600 2887.4100 3055.2600 2889.4100 ;
        RECT 3292.7200 2887.4100 3295.7200 2889.4100 ;
        RECT 3533.1800 2637.5700 3536.1800 2639.5700 ;
        RECT 3783.0700 2638.5700 3784.5700 2640.0700 ;
        RECT 3533.1800 2887.4100 3536.1800 2889.4100 ;
        RECT 3783.0700 2888.4100 3784.5700 2889.9100 ;
        RECT 2090.4200 3137.2500 2093.4200 3139.2500 ;
        RECT 2330.8800 3137.2500 2333.8800 3139.2500 ;
        RECT 2090.4200 3387.0900 2093.4200 3389.0900 ;
        RECT 2330.8800 3387.0900 2333.8800 3389.0900 ;
        RECT 2571.3400 3137.2500 2574.3400 3139.2500 ;
        RECT 2811.8000 3137.2500 2814.8000 3139.2500 ;
        RECT 2571.3400 3387.0900 2574.3400 3389.0900 ;
        RECT 2811.8000 3387.0900 2814.8000 3389.0900 ;
        RECT 2090.4200 3636.9300 2093.4200 3638.9300 ;
        RECT 2330.8800 3636.9300 2333.8800 3638.9300 ;
        RECT 2091.4200 3910.8400 2093.4200 3912.8400 ;
        RECT 2331.8800 3910.8400 2333.8800 3912.8400 ;
        RECT 2811.8000 3636.9300 2814.8000 3638.9300 ;
        RECT 2572.3400 3910.8400 2574.3400 3912.8400 ;
        RECT 2812.8000 3910.8400 2814.8000 3912.8400 ;
        RECT 3052.2600 3137.2500 3055.2600 3139.2500 ;
        RECT 3292.7200 3137.2500 3295.7200 3139.2500 ;
        RECT 3052.2600 3387.0900 3055.2600 3389.0900 ;
        RECT 3292.7200 3387.0900 3295.7200 3389.0900 ;
        RECT 3533.1800 3137.2500 3536.1800 3139.2500 ;
        RECT 3783.0700 3138.2500 3784.5700 3139.7500 ;
        RECT 3533.1800 3387.0900 3536.1800 3389.0900 ;
        RECT 3783.0700 3388.0900 3784.5700 3389.5900 ;
        RECT 3052.2600 3636.9300 3055.2600 3638.9300 ;
        RECT 3292.7200 3636.9300 3295.7200 3638.9300 ;
        RECT 3053.2600 3910.8400 3055.2600 3912.8400 ;
        RECT 3293.7200 3910.8400 3295.7200 3912.8400 ;
        RECT 3533.1800 3636.9300 3536.1800 3638.9300 ;
        RECT 3783.0700 3637.9300 3784.5700 3639.4300 ;
        RECT 3534.1800 3910.8400 3536.1800 3912.8400 ;
        RECT 153.3400 140.4300 156.0100 141.9300 ;
        RECT 153.3400 390.2700 156.0100 391.7700 ;
        RECT 153.3400 640.1100 156.0100 641.6100 ;
        RECT 153.3400 889.9500 156.0100 891.4500 ;
        RECT 153.3400 1139.7900 156.0100 1141.2900 ;
        RECT 153.3400 1389.6300 156.0100 1391.1300 ;
        RECT 153.3400 1639.4700 156.0100 1640.9700 ;
        RECT 153.3400 1889.3100 156.0100 1890.8100 ;
        RECT 153.3400 2139.1500 156.0100 2140.6500 ;
        RECT 153.3400 2388.9900 156.0100 2390.4900 ;
        RECT 153.3400 2638.8300 156.0100 2640.3300 ;
        RECT 153.3400 2888.6700 156.0100 2890.1700 ;
        RECT 153.3400 3138.5100 156.0100 3140.0100 ;
        RECT 153.3400 3388.3500 156.0100 3389.8500 ;
        RECT 153.3400 3638.1900 156.0100 3639.6900 ;
      LAYER met5 ;
        RECT 161.0800 129.2400 3819.9800 131.2400 ;
        RECT 8.0000 78.9800 3770.0800 80.9800 ;
        RECT 8.0000 8.0000 3922.2400 12.0000 ;
        RECT 161.0800 379.0800 3819.9800 381.0800 ;
        RECT 161.0800 628.9200 3819.9800 630.9200 ;
        RECT 161.0800 878.7600 3819.9800 880.7600 ;
        RECT 161.0800 1878.1200 3819.9800 1880.1200 ;
        RECT 161.0800 1628.2800 3819.9800 1630.2800 ;
        RECT 161.0800 1378.4400 3819.9800 1380.4400 ;
        RECT 161.0800 1128.6000 3819.9800 1130.6000 ;
        RECT 8.0000 129.5000 163.0800 131.5000 ;
        RECT 153.3400 140.3800 163.0800 141.9800 ;
        RECT 117.1800 373.3400 163.0800 375.3400 ;
        RECT 8.0000 379.3400 163.0800 381.3400 ;
        RECT 153.3400 390.2200 163.0800 391.8200 ;
        RECT 8.0000 629.1800 163.0800 631.1800 ;
        RECT 117.1800 623.1800 163.0800 625.1800 ;
        RECT 153.3400 640.0600 163.0800 641.6600 ;
        RECT 117.1800 873.0200 163.0800 875.0200 ;
        RECT 8.0000 879.0200 163.0800 881.0200 ;
        RECT 153.3400 889.9000 163.0800 891.5000 ;
        RECT 117.1800 1122.8600 163.0800 1124.8600 ;
        RECT 8.0000 1128.8600 163.0800 1130.8600 ;
        RECT 153.3400 1139.7400 163.0800 1141.3400 ;
        RECT 117.1800 1372.7000 163.0800 1374.7000 ;
        RECT 8.0000 1378.7000 163.0800 1380.7000 ;
        RECT 153.3400 1389.5800 163.0800 1391.1800 ;
        RECT 117.1800 1622.5400 163.0800 1624.5400 ;
        RECT 8.0000 1628.5400 163.0800 1630.5400 ;
        RECT 153.3400 1639.4200 163.0800 1641.0200 ;
        RECT 117.1800 1872.3800 163.0800 1874.3800 ;
        RECT 8.0000 1878.3800 163.0800 1880.3800 ;
        RECT 153.3400 1889.2600 163.0800 1890.8600 ;
        RECT 8.0000 3918.0600 3922.2400 3922.0600 ;
        RECT 161.0800 2127.9600 3819.9800 2129.9600 ;
        RECT 161.0800 2377.8000 3819.9800 2379.8000 ;
        RECT 161.0800 2627.6400 3819.9800 2629.6400 ;
        RECT 161.0800 2877.4800 3819.9800 2879.4800 ;
        RECT 161.0800 3127.3200 3819.9800 3129.3200 ;
        RECT 161.0800 3377.1600 3819.9800 3379.1600 ;
        RECT 161.0800 3627.0000 3819.9800 3629.0000 ;
        RECT 161.0800 3876.8400 3770.0800 3878.8400 ;
        RECT 117.1800 2122.2200 163.0800 2124.2200 ;
        RECT 8.0000 2128.2200 163.0800 2130.2200 ;
        RECT 153.3400 2139.1000 163.0800 2140.7000 ;
        RECT 8.0000 2378.0600 163.0800 2380.0600 ;
        RECT 117.1800 2372.0600 163.0800 2374.0600 ;
        RECT 153.3400 2388.9400 163.0800 2390.5400 ;
        RECT 117.1800 2621.9000 163.0800 2623.9000 ;
        RECT 8.0000 2627.9000 163.0800 2629.9000 ;
        RECT 153.3400 2638.7800 163.0800 2640.3800 ;
        RECT 117.1800 2871.7400 163.0800 2873.7400 ;
        RECT 8.0000 2877.7400 163.0800 2879.7400 ;
        RECT 153.3400 2888.6200 163.0800 2890.2200 ;
        RECT 117.1800 3121.5800 163.0800 3123.5800 ;
        RECT 8.0000 3127.5800 163.0800 3129.5800 ;
        RECT 153.3400 3138.4600 163.0800 3140.0600 ;
        RECT 8.0000 3377.4200 163.0800 3379.4200 ;
        RECT 117.1800 3371.4200 163.0800 3373.4200 ;
        RECT 153.3400 3388.3000 163.0800 3389.9000 ;
        RECT 117.1800 3621.2600 163.0800 3623.2600 ;
        RECT 8.0000 3627.2600 163.0800 3629.2600 ;
        RECT 153.3400 3638.1400 163.0800 3639.7400 ;
        RECT 8.0000 3871.1000 163.0800 3873.1000 ;
        RECT 161.0800 140.1800 163.0800 142.1800 ;
        RECT 161.0800 129.2400 163.0800 131.5000 ;
        RECT 161.0800 379.0800 163.0800 381.3400 ;
        RECT 161.0800 390.0200 163.0800 392.0200 ;
        RECT 161.0800 628.9200 163.0800 631.1800 ;
        RECT 161.0800 639.8600 163.0800 641.8600 ;
        RECT 161.0800 878.7600 163.0800 881.0200 ;
        RECT 161.0800 889.7000 163.0800 891.7000 ;
        RECT 161.0800 1128.6000 163.0800 1130.8600 ;
        RECT 161.0800 1139.5400 163.0800 1141.5400 ;
        RECT 161.0800 1378.4400 163.0800 1380.7000 ;
        RECT 161.0800 1389.3800 163.0800 1391.3800 ;
        RECT 161.0800 1628.2800 163.0800 1630.5400 ;
        RECT 161.0800 1639.2200 163.0800 1641.2200 ;
        RECT 161.0800 1878.1200 163.0800 1880.3800 ;
        RECT 161.0800 1889.0600 163.0800 1891.0600 ;
        RECT 161.0800 2127.9600 163.0800 2130.2200 ;
        RECT 161.0800 2138.9000 163.0800 2140.9000 ;
        RECT 161.0800 2377.8000 163.0800 2380.0600 ;
        RECT 161.0800 2388.7400 163.0800 2390.7400 ;
        RECT 161.0800 2627.6400 163.0800 2629.9000 ;
        RECT 161.0800 2638.5800 163.0800 2640.5800 ;
        RECT 161.0800 2877.4800 163.0800 2879.7400 ;
        RECT 161.0800 2888.4200 163.0800 2890.4200 ;
        RECT 161.0800 3127.3200 163.0800 3129.5800 ;
        RECT 161.0800 3138.2600 163.0800 3140.2600 ;
        RECT 161.0800 3377.1600 163.0800 3379.4200 ;
        RECT 161.0800 3388.1000 163.0800 3390.1000 ;
        RECT 161.0800 3627.0000 163.0800 3629.2600 ;
        RECT 161.0800 3637.9400 163.0800 3639.9400 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 3930.2400 3930.0600 ;
    LAYER met1 ;
      RECT 0.0000 3745.4800 3930.2400 3930.0600 ;
      RECT 0.7350 3745.1400 3930.2400 3745.4800 ;
      RECT 0.7350 3745.0600 3929.5050 3745.1400 ;
      RECT 0.0000 3744.7200 3929.5050 3745.0600 ;
      RECT 0.0000 3743.4400 3930.2400 3744.7200 ;
      RECT 0.0000 3743.0200 3929.5050 3743.4400 ;
      RECT 0.0000 3741.7400 3930.2400 3743.0200 ;
      RECT 0.0000 3741.4000 3929.5050 3741.7400 ;
      RECT 0.7350 3741.3200 3929.5050 3741.4000 ;
      RECT 0.7350 3740.9800 3930.2400 3741.3200 ;
      RECT 0.0000 3740.3800 3930.2400 3740.9800 ;
      RECT 0.0000 3739.9600 3929.5050 3740.3800 ;
      RECT 0.0000 3738.6800 3930.2400 3739.9600 ;
      RECT 0.0000 3738.2600 3929.5050 3738.6800 ;
      RECT 0.0000 3737.3200 3930.2400 3738.2600 ;
      RECT 0.7350 3736.9800 3930.2400 3737.3200 ;
      RECT 0.7350 3736.9000 3929.5050 3736.9800 ;
      RECT 0.0000 3736.5600 3929.5050 3736.9000 ;
      RECT 0.0000 3735.6200 3930.2400 3736.5600 ;
      RECT 0.0000 3735.2000 3929.5050 3735.6200 ;
      RECT 0.0000 3733.9200 3930.2400 3735.2000 ;
      RECT 0.0000 3733.5800 3929.5050 3733.9200 ;
      RECT 0.7350 3733.5000 3929.5050 3733.5800 ;
      RECT 0.7350 3733.1600 3930.2400 3733.5000 ;
      RECT 0.0000 3732.2200 3930.2400 3733.1600 ;
      RECT 0.0000 3731.8000 3929.5050 3732.2200 ;
      RECT 0.0000 3730.8600 3930.2400 3731.8000 ;
      RECT 0.0000 3730.4400 3929.5050 3730.8600 ;
      RECT 0.0000 3729.5000 3930.2400 3730.4400 ;
      RECT 0.7350 3729.1600 3930.2400 3729.5000 ;
      RECT 0.7350 3729.0800 3929.5050 3729.1600 ;
      RECT 0.0000 3728.7400 3929.5050 3729.0800 ;
      RECT 0.0000 3727.8000 3930.2400 3728.7400 ;
      RECT 0.0000 3727.3800 3929.5050 3727.8000 ;
      RECT 0.0000 3726.1000 3930.2400 3727.3800 ;
      RECT 0.0000 3725.7600 3929.5050 3726.1000 ;
      RECT 0.7350 3725.6800 3929.5050 3725.7600 ;
      RECT 0.7350 3725.3400 3930.2400 3725.6800 ;
      RECT 0.0000 3724.4000 3930.2400 3725.3400 ;
      RECT 0.0000 3723.9800 3929.5050 3724.4000 ;
      RECT 0.0000 3723.0400 3930.2400 3723.9800 ;
      RECT 0.0000 3722.6200 3929.5050 3723.0400 ;
      RECT 0.0000 3721.3400 3930.2400 3722.6200 ;
      RECT 0.0000 3720.9200 3929.5050 3721.3400 ;
      RECT 0.0000 3719.6400 3930.2400 3720.9200 ;
      RECT 0.0000 3719.2200 3929.5050 3719.6400 ;
      RECT 0.0000 3718.2800 3930.2400 3719.2200 ;
      RECT 0.0000 3717.8600 3929.5050 3718.2800 ;
      RECT 0.0000 3716.5800 3930.2400 3717.8600 ;
      RECT 0.0000 3716.1600 3929.5050 3716.5800 ;
      RECT 0.0000 3715.2200 3930.2400 3716.1600 ;
      RECT 0.0000 3714.8000 3929.5050 3715.2200 ;
      RECT 0.0000 3495.5800 3930.2400 3714.8000 ;
      RECT 0.7350 3495.2400 3930.2400 3495.5800 ;
      RECT 0.7350 3495.1600 3929.5050 3495.2400 ;
      RECT 0.0000 3494.8200 3929.5050 3495.1600 ;
      RECT 0.0000 3493.5400 3930.2400 3494.8200 ;
      RECT 0.0000 3493.1200 3929.5050 3493.5400 ;
      RECT 0.0000 3491.8400 3930.2400 3493.1200 ;
      RECT 0.0000 3491.5000 3929.5050 3491.8400 ;
      RECT 0.7350 3491.4200 3929.5050 3491.5000 ;
      RECT 0.7350 3491.0800 3930.2400 3491.4200 ;
      RECT 0.0000 3490.4800 3930.2400 3491.0800 ;
      RECT 0.0000 3490.0600 3929.5050 3490.4800 ;
      RECT 0.0000 3488.7800 3930.2400 3490.0600 ;
      RECT 0.0000 3488.3600 3929.5050 3488.7800 ;
      RECT 0.0000 3487.4200 3930.2400 3488.3600 ;
      RECT 0.7350 3487.0800 3930.2400 3487.4200 ;
      RECT 0.7350 3487.0000 3929.5050 3487.0800 ;
      RECT 0.0000 3486.6600 3929.5050 3487.0000 ;
      RECT 0.0000 3485.7200 3930.2400 3486.6600 ;
      RECT 0.0000 3485.3000 3929.5050 3485.7200 ;
      RECT 0.0000 3484.0200 3930.2400 3485.3000 ;
      RECT 0.0000 3483.6800 3929.5050 3484.0200 ;
      RECT 0.7350 3483.6000 3929.5050 3483.6800 ;
      RECT 0.7350 3483.2600 3930.2400 3483.6000 ;
      RECT 0.0000 3482.3200 3930.2400 3483.2600 ;
      RECT 0.0000 3481.9000 3929.5050 3482.3200 ;
      RECT 0.0000 3480.9600 3930.2400 3481.9000 ;
      RECT 0.0000 3480.5400 3929.5050 3480.9600 ;
      RECT 0.0000 3479.6000 3930.2400 3480.5400 ;
      RECT 0.7350 3479.2600 3930.2400 3479.6000 ;
      RECT 0.7350 3479.1800 3929.5050 3479.2600 ;
      RECT 0.0000 3478.8400 3929.5050 3479.1800 ;
      RECT 0.0000 3477.9000 3930.2400 3478.8400 ;
      RECT 0.0000 3477.4800 3929.5050 3477.9000 ;
      RECT 0.0000 3476.2000 3930.2400 3477.4800 ;
      RECT 0.0000 3475.8600 3929.5050 3476.2000 ;
      RECT 0.7350 3475.7800 3929.5050 3475.8600 ;
      RECT 0.7350 3475.4400 3930.2400 3475.7800 ;
      RECT 0.0000 3474.5000 3930.2400 3475.4400 ;
      RECT 0.0000 3474.0800 3929.5050 3474.5000 ;
      RECT 0.0000 3473.1400 3930.2400 3474.0800 ;
      RECT 0.0000 3472.7200 3929.5050 3473.1400 ;
      RECT 0.0000 3471.4400 3930.2400 3472.7200 ;
      RECT 0.0000 3471.0200 3929.5050 3471.4400 ;
      RECT 0.0000 3469.7400 3930.2400 3471.0200 ;
      RECT 0.0000 3469.3200 3929.5050 3469.7400 ;
      RECT 0.0000 3468.7200 3930.2400 3469.3200 ;
      RECT 0.0000 3468.3000 3929.5050 3468.7200 ;
      RECT 0.0000 3466.6800 3930.2400 3468.3000 ;
      RECT 0.0000 3466.2600 3929.5050 3466.6800 ;
      RECT 0.0000 3465.6600 3930.2400 3466.2600 ;
      RECT 0.0000 3465.2400 3929.5050 3465.6600 ;
      RECT 0.0000 3245.6800 3930.2400 3465.2400 ;
      RECT 0.7350 3245.2600 3929.5050 3245.6800 ;
      RECT 0.0000 3243.9800 3930.2400 3245.2600 ;
      RECT 0.0000 3243.5600 3929.5050 3243.9800 ;
      RECT 0.0000 3242.2800 3930.2400 3243.5600 ;
      RECT 0.0000 3241.8600 3929.5050 3242.2800 ;
      RECT 0.0000 3241.6000 3930.2400 3241.8600 ;
      RECT 0.7350 3241.1800 3930.2400 3241.6000 ;
      RECT 0.0000 3240.9200 3930.2400 3241.1800 ;
      RECT 0.0000 3240.5000 3929.5050 3240.9200 ;
      RECT 0.0000 3239.2200 3930.2400 3240.5000 ;
      RECT 0.0000 3238.8000 3929.5050 3239.2200 ;
      RECT 0.0000 3237.5200 3930.2400 3238.8000 ;
      RECT 0.7350 3237.1000 3929.5050 3237.5200 ;
      RECT 0.0000 3236.1600 3930.2400 3237.1000 ;
      RECT 0.0000 3235.7400 3929.5050 3236.1600 ;
      RECT 0.0000 3234.4600 3930.2400 3235.7400 ;
      RECT 0.0000 3234.0400 3929.5050 3234.4600 ;
      RECT 0.0000 3233.7800 3930.2400 3234.0400 ;
      RECT 0.7350 3233.3600 3930.2400 3233.7800 ;
      RECT 0.0000 3232.4200 3930.2400 3233.3600 ;
      RECT 0.0000 3232.0000 3929.5050 3232.4200 ;
      RECT 0.0000 3231.4000 3930.2400 3232.0000 ;
      RECT 0.0000 3230.9800 3929.5050 3231.4000 ;
      RECT 0.0000 3229.7000 3930.2400 3230.9800 ;
      RECT 0.7350 3229.3600 3930.2400 3229.7000 ;
      RECT 0.7350 3229.2800 3929.5050 3229.3600 ;
      RECT 0.0000 3228.9400 3929.5050 3229.2800 ;
      RECT 0.0000 3228.3400 3930.2400 3228.9400 ;
      RECT 0.0000 3227.9200 3929.5050 3228.3400 ;
      RECT 0.0000 3226.3000 3930.2400 3227.9200 ;
      RECT 0.0000 3225.9600 3929.5050 3226.3000 ;
      RECT 0.7350 3225.8800 3929.5050 3225.9600 ;
      RECT 0.7350 3225.5400 3930.2400 3225.8800 ;
      RECT 0.0000 3224.9400 3930.2400 3225.5400 ;
      RECT 0.0000 3224.5200 3929.5050 3224.9400 ;
      RECT 0.0000 3223.2400 3930.2400 3224.5200 ;
      RECT 0.0000 3222.8200 3929.5050 3223.2400 ;
      RECT 0.0000 3221.8800 3930.2400 3222.8200 ;
      RECT 0.0000 3221.4600 3929.5050 3221.8800 ;
      RECT 0.0000 3220.1800 3930.2400 3221.4600 ;
      RECT 0.0000 3219.7600 3929.5050 3220.1800 ;
      RECT 0.0000 3218.8200 3930.2400 3219.7600 ;
      RECT 0.0000 3218.4000 3929.5050 3218.8200 ;
      RECT 0.0000 3217.1200 3930.2400 3218.4000 ;
      RECT 0.0000 3216.7000 3929.5050 3217.1200 ;
      RECT 0.0000 3215.7600 3930.2400 3216.7000 ;
      RECT 0.0000 3215.3400 3929.5050 3215.7600 ;
      RECT 0.0000 2995.7800 3930.2400 3215.3400 ;
      RECT 0.7350 2995.3600 3929.5050 2995.7800 ;
      RECT 0.0000 2994.0800 3930.2400 2995.3600 ;
      RECT 0.0000 2993.6600 3929.5050 2994.0800 ;
      RECT 0.0000 2992.3800 3930.2400 2993.6600 ;
      RECT 0.0000 2991.9600 3929.5050 2992.3800 ;
      RECT 0.0000 2991.7000 3930.2400 2991.9600 ;
      RECT 0.7350 2991.2800 3930.2400 2991.7000 ;
      RECT 0.0000 2991.0200 3930.2400 2991.2800 ;
      RECT 0.0000 2990.6000 3929.5050 2991.0200 ;
      RECT 0.0000 2989.3200 3930.2400 2990.6000 ;
      RECT 0.0000 2988.9000 3929.5050 2989.3200 ;
      RECT 0.0000 2987.9600 3930.2400 2988.9000 ;
      RECT 0.7350 2987.6200 3930.2400 2987.9600 ;
      RECT 0.7350 2987.5400 3929.5050 2987.6200 ;
      RECT 0.0000 2987.2000 3929.5050 2987.5400 ;
      RECT 0.0000 2986.2600 3930.2400 2987.2000 ;
      RECT 0.0000 2985.8400 3929.5050 2986.2600 ;
      RECT 0.0000 2984.5600 3930.2400 2985.8400 ;
      RECT 0.0000 2984.1400 3929.5050 2984.5600 ;
      RECT 0.0000 2983.8800 3930.2400 2984.1400 ;
      RECT 0.7350 2983.4600 3930.2400 2983.8800 ;
      RECT 0.0000 2982.8600 3930.2400 2983.4600 ;
      RECT 0.0000 2982.4400 3929.5050 2982.8600 ;
      RECT 0.0000 2981.5000 3930.2400 2982.4400 ;
      RECT 0.0000 2981.0800 3929.5050 2981.5000 ;
      RECT 0.0000 2979.8000 3930.2400 2981.0800 ;
      RECT 0.7350 2979.3800 3929.5050 2979.8000 ;
      RECT 0.0000 2978.4400 3930.2400 2979.3800 ;
      RECT 0.0000 2978.0200 3929.5050 2978.4400 ;
      RECT 0.0000 2976.7400 3930.2400 2978.0200 ;
      RECT 0.0000 2976.4000 3929.5050 2976.7400 ;
      RECT 0.7350 2976.3200 3929.5050 2976.4000 ;
      RECT 0.7350 2975.9800 3930.2400 2976.3200 ;
      RECT 0.0000 2975.0400 3930.2400 2975.9800 ;
      RECT 0.0000 2974.6200 3929.5050 2975.0400 ;
      RECT 0.0000 2973.6800 3930.2400 2974.6200 ;
      RECT 0.0000 2973.2600 3929.5050 2973.6800 ;
      RECT 0.0000 2971.9800 3930.2400 2973.2600 ;
      RECT 0.0000 2971.5600 3929.5050 2971.9800 ;
      RECT 0.0000 2970.2800 3930.2400 2971.5600 ;
      RECT 0.0000 2969.8600 3929.5050 2970.2800 ;
      RECT 0.0000 2968.9200 3930.2400 2969.8600 ;
      RECT 0.0000 2968.5000 3929.5050 2968.9200 ;
      RECT 0.0000 2967.2200 3930.2400 2968.5000 ;
      RECT 0.0000 2966.8000 3929.5050 2967.2200 ;
      RECT 0.0000 2965.8600 3930.2400 2966.8000 ;
      RECT 0.0000 2965.4400 3929.5050 2965.8600 ;
      RECT 0.0000 2746.2200 3930.2400 2965.4400 ;
      RECT 0.7350 2745.8800 3930.2400 2746.2200 ;
      RECT 0.7350 2745.8000 3929.5050 2745.8800 ;
      RECT 0.0000 2745.4600 3929.5050 2745.8000 ;
      RECT 0.0000 2744.1800 3930.2400 2745.4600 ;
      RECT 0.0000 2743.7600 3929.5050 2744.1800 ;
      RECT 0.0000 2742.4800 3930.2400 2743.7600 ;
      RECT 0.0000 2742.1400 3929.5050 2742.4800 ;
      RECT 0.7350 2742.0600 3929.5050 2742.1400 ;
      RECT 0.7350 2741.7200 3930.2400 2742.0600 ;
      RECT 0.0000 2741.1200 3930.2400 2741.7200 ;
      RECT 0.0000 2740.7000 3929.5050 2741.1200 ;
      RECT 0.0000 2739.4200 3930.2400 2740.7000 ;
      RECT 0.0000 2739.0000 3929.5050 2739.4200 ;
      RECT 0.0000 2738.0600 3930.2400 2739.0000 ;
      RECT 0.7350 2737.7200 3930.2400 2738.0600 ;
      RECT 0.7350 2737.6400 3929.5050 2737.7200 ;
      RECT 0.0000 2737.3000 3929.5050 2737.6400 ;
      RECT 0.0000 2736.3600 3930.2400 2737.3000 ;
      RECT 0.0000 2735.9400 3929.5050 2736.3600 ;
      RECT 0.0000 2734.6600 3930.2400 2735.9400 ;
      RECT 0.0000 2734.2400 3929.5050 2734.6600 ;
      RECT 0.0000 2733.9800 3930.2400 2734.2400 ;
      RECT 0.7350 2733.5600 3930.2400 2733.9800 ;
      RECT 0.0000 2732.9600 3930.2400 2733.5600 ;
      RECT 0.0000 2732.5400 3929.5050 2732.9600 ;
      RECT 0.0000 2731.6000 3930.2400 2732.5400 ;
      RECT 0.0000 2731.1800 3929.5050 2731.6000 ;
      RECT 0.0000 2730.2400 3930.2400 2731.1800 ;
      RECT 0.7350 2729.9000 3930.2400 2730.2400 ;
      RECT 0.7350 2729.8200 3929.5050 2729.9000 ;
      RECT 0.0000 2729.4800 3929.5050 2729.8200 ;
      RECT 0.0000 2728.5400 3930.2400 2729.4800 ;
      RECT 0.0000 2728.1200 3929.5050 2728.5400 ;
      RECT 0.0000 2726.8400 3930.2400 2728.1200 ;
      RECT 0.0000 2726.5000 3929.5050 2726.8400 ;
      RECT 0.7350 2726.4200 3929.5050 2726.5000 ;
      RECT 0.7350 2726.0800 3930.2400 2726.4200 ;
      RECT 0.0000 2725.1400 3930.2400 2726.0800 ;
      RECT 0.0000 2724.7200 3929.5050 2725.1400 ;
      RECT 0.0000 2723.7800 3930.2400 2724.7200 ;
      RECT 0.0000 2723.3600 3929.5050 2723.7800 ;
      RECT 0.0000 2722.0800 3930.2400 2723.3600 ;
      RECT 0.0000 2721.6600 3929.5050 2722.0800 ;
      RECT 0.0000 2720.3800 3930.2400 2721.6600 ;
      RECT 0.0000 2719.9600 3929.5050 2720.3800 ;
      RECT 0.0000 2719.0200 3930.2400 2719.9600 ;
      RECT 0.0000 2718.6000 3929.5050 2719.0200 ;
      RECT 0.0000 2717.3200 3930.2400 2718.6000 ;
      RECT 0.0000 2716.9000 3929.5050 2717.3200 ;
      RECT 0.0000 2715.9600 3930.2400 2716.9000 ;
      RECT 0.0000 2715.5400 3929.5050 2715.9600 ;
      RECT 0.0000 2496.3200 3930.2400 2715.5400 ;
      RECT 0.7350 2495.9800 3930.2400 2496.3200 ;
      RECT 0.7350 2495.9000 3929.5050 2495.9800 ;
      RECT 0.0000 2495.5600 3929.5050 2495.9000 ;
      RECT 0.0000 2494.2800 3930.2400 2495.5600 ;
      RECT 0.0000 2493.8600 3929.5050 2494.2800 ;
      RECT 0.0000 2492.5800 3930.2400 2493.8600 ;
      RECT 0.0000 2492.2400 3929.5050 2492.5800 ;
      RECT 0.7350 2492.1600 3929.5050 2492.2400 ;
      RECT 0.7350 2491.8200 3930.2400 2492.1600 ;
      RECT 0.0000 2491.2200 3930.2400 2491.8200 ;
      RECT 0.0000 2490.8000 3929.5050 2491.2200 ;
      RECT 0.0000 2489.5200 3930.2400 2490.8000 ;
      RECT 0.0000 2489.1000 3929.5050 2489.5200 ;
      RECT 0.0000 2488.1600 3930.2400 2489.1000 ;
      RECT 0.7350 2487.8200 3930.2400 2488.1600 ;
      RECT 0.7350 2487.7400 3929.5050 2487.8200 ;
      RECT 0.0000 2487.4000 3929.5050 2487.7400 ;
      RECT 0.0000 2486.4600 3930.2400 2487.4000 ;
      RECT 0.0000 2486.0400 3929.5050 2486.4600 ;
      RECT 0.0000 2484.7600 3930.2400 2486.0400 ;
      RECT 0.0000 2484.4200 3929.5050 2484.7600 ;
      RECT 0.7350 2484.3400 3929.5050 2484.4200 ;
      RECT 0.7350 2484.0000 3930.2400 2484.3400 ;
      RECT 0.0000 2483.0600 3930.2400 2484.0000 ;
      RECT 0.0000 2482.6400 3929.5050 2483.0600 ;
      RECT 0.0000 2481.7000 3930.2400 2482.6400 ;
      RECT 0.0000 2481.2800 3929.5050 2481.7000 ;
      RECT 0.0000 2480.3400 3930.2400 2481.2800 ;
      RECT 0.7350 2480.0000 3930.2400 2480.3400 ;
      RECT 0.7350 2479.9200 3929.5050 2480.0000 ;
      RECT 0.0000 2479.5800 3929.5050 2479.9200 ;
      RECT 0.0000 2478.6400 3930.2400 2479.5800 ;
      RECT 0.0000 2478.2200 3929.5050 2478.6400 ;
      RECT 0.0000 2476.9400 3930.2400 2478.2200 ;
      RECT 0.0000 2476.6000 3929.5050 2476.9400 ;
      RECT 0.7350 2476.5200 3929.5050 2476.6000 ;
      RECT 0.7350 2476.1800 3930.2400 2476.5200 ;
      RECT 0.0000 2475.2400 3930.2400 2476.1800 ;
      RECT 0.0000 2474.8200 3929.5050 2475.2400 ;
      RECT 0.0000 2473.8800 3930.2400 2474.8200 ;
      RECT 0.0000 2473.4600 3929.5050 2473.8800 ;
      RECT 0.0000 2472.1800 3930.2400 2473.4600 ;
      RECT 0.0000 2471.7600 3929.5050 2472.1800 ;
      RECT 0.0000 2470.4800 3930.2400 2471.7600 ;
      RECT 0.0000 2470.0600 3929.5050 2470.4800 ;
      RECT 0.0000 2469.1200 3930.2400 2470.0600 ;
      RECT 0.0000 2468.7000 3929.5050 2469.1200 ;
      RECT 0.0000 2467.4200 3930.2400 2468.7000 ;
      RECT 0.0000 2467.0000 3929.5050 2467.4200 ;
      RECT 0.0000 2466.0600 3930.2400 2467.0000 ;
      RECT 0.0000 2465.6400 3929.5050 2466.0600 ;
      RECT 0.0000 2246.4200 3930.2400 2465.6400 ;
      RECT 0.7350 2246.0800 3930.2400 2246.4200 ;
      RECT 0.7350 2246.0000 3929.5050 2246.0800 ;
      RECT 0.0000 2245.6600 3929.5050 2246.0000 ;
      RECT 0.0000 2244.3800 3930.2400 2245.6600 ;
      RECT 0.0000 2243.9600 3929.5050 2244.3800 ;
      RECT 0.0000 2242.6800 3930.2400 2243.9600 ;
      RECT 0.0000 2242.3400 3929.5050 2242.6800 ;
      RECT 0.7350 2242.2600 3929.5050 2242.3400 ;
      RECT 0.7350 2241.9200 3930.2400 2242.2600 ;
      RECT 0.0000 2241.3200 3930.2400 2241.9200 ;
      RECT 0.0000 2240.9000 3929.5050 2241.3200 ;
      RECT 0.0000 2239.6200 3930.2400 2240.9000 ;
      RECT 0.0000 2239.2000 3929.5050 2239.6200 ;
      RECT 0.0000 2238.2600 3930.2400 2239.2000 ;
      RECT 0.7350 2237.9200 3930.2400 2238.2600 ;
      RECT 0.7350 2237.8400 3929.5050 2237.9200 ;
      RECT 0.0000 2237.5000 3929.5050 2237.8400 ;
      RECT 0.0000 2236.5600 3930.2400 2237.5000 ;
      RECT 0.0000 2236.1400 3929.5050 2236.5600 ;
      RECT 0.0000 2234.8600 3930.2400 2236.1400 ;
      RECT 0.0000 2234.5200 3929.5050 2234.8600 ;
      RECT 0.7350 2234.4400 3929.5050 2234.5200 ;
      RECT 0.7350 2234.1000 3930.2400 2234.4400 ;
      RECT 0.0000 2233.1600 3930.2400 2234.1000 ;
      RECT 0.0000 2232.7400 3929.5050 2233.1600 ;
      RECT 0.0000 2231.8000 3930.2400 2232.7400 ;
      RECT 0.0000 2231.3800 3929.5050 2231.8000 ;
      RECT 0.0000 2230.4400 3930.2400 2231.3800 ;
      RECT 0.7350 2230.1000 3930.2400 2230.4400 ;
      RECT 0.7350 2230.0200 3929.5050 2230.1000 ;
      RECT 0.0000 2229.6800 3929.5050 2230.0200 ;
      RECT 0.0000 2228.7400 3930.2400 2229.6800 ;
      RECT 0.0000 2228.3200 3929.5050 2228.7400 ;
      RECT 0.0000 2227.0400 3930.2400 2228.3200 ;
      RECT 0.0000 2226.7000 3929.5050 2227.0400 ;
      RECT 0.7350 2226.6200 3929.5050 2226.7000 ;
      RECT 0.7350 2226.2800 3930.2400 2226.6200 ;
      RECT 0.0000 2225.3400 3930.2400 2226.2800 ;
      RECT 0.0000 2224.9200 3929.5050 2225.3400 ;
      RECT 0.0000 2223.9800 3930.2400 2224.9200 ;
      RECT 0.0000 2223.5600 3929.5050 2223.9800 ;
      RECT 0.0000 2222.2800 3930.2400 2223.5600 ;
      RECT 0.0000 2221.8600 3929.5050 2222.2800 ;
      RECT 0.0000 2220.5800 3930.2400 2221.8600 ;
      RECT 0.0000 2220.1600 3929.5050 2220.5800 ;
      RECT 0.0000 2219.2200 3930.2400 2220.1600 ;
      RECT 0.0000 2218.8000 3929.5050 2219.2200 ;
      RECT 0.0000 2217.5200 3930.2400 2218.8000 ;
      RECT 0.0000 2217.1000 3929.5050 2217.5200 ;
      RECT 0.0000 2216.1600 3930.2400 2217.1000 ;
      RECT 0.0000 2215.7400 3929.5050 2216.1600 ;
      RECT 0.0000 1996.5200 3930.2400 2215.7400 ;
      RECT 0.7350 1996.1800 3930.2400 1996.5200 ;
      RECT 0.7350 1996.1000 3929.5050 1996.1800 ;
      RECT 0.0000 1995.7600 3929.5050 1996.1000 ;
      RECT 0.0000 1994.4800 3930.2400 1995.7600 ;
      RECT 0.0000 1994.0600 3929.5050 1994.4800 ;
      RECT 0.0000 1993.1200 3930.2400 1994.0600 ;
      RECT 0.0000 1992.7000 3929.5050 1993.1200 ;
      RECT 0.0000 1992.4400 3930.2400 1992.7000 ;
      RECT 0.7350 1992.0200 3930.2400 1992.4400 ;
      RECT 0.0000 1991.4200 3930.2400 1992.0200 ;
      RECT 0.0000 1991.0000 3929.5050 1991.4200 ;
      RECT 0.0000 1990.0600 3930.2400 1991.0000 ;
      RECT 0.0000 1989.6400 3929.5050 1990.0600 ;
      RECT 0.0000 1988.3600 3930.2400 1989.6400 ;
      RECT 0.7350 1988.0200 3930.2400 1988.3600 ;
      RECT 0.7350 1987.9400 3929.5050 1988.0200 ;
      RECT 0.0000 1987.6000 3929.5050 1987.9400 ;
      RECT 0.0000 1987.0000 3930.2400 1987.6000 ;
      RECT 0.0000 1986.5800 3929.5050 1987.0000 ;
      RECT 0.0000 1984.9600 3930.2400 1986.5800 ;
      RECT 0.0000 1984.6200 3929.5050 1984.9600 ;
      RECT 0.7350 1984.5400 3929.5050 1984.6200 ;
      RECT 0.7350 1984.2000 3930.2400 1984.5400 ;
      RECT 0.0000 1983.2600 3930.2400 1984.2000 ;
      RECT 0.0000 1982.8400 3929.5050 1983.2600 ;
      RECT 0.0000 1981.9000 3930.2400 1982.8400 ;
      RECT 0.0000 1981.4800 3929.5050 1981.9000 ;
      RECT 0.0000 1980.5400 3930.2400 1981.4800 ;
      RECT 0.7350 1980.2000 3930.2400 1980.5400 ;
      RECT 0.7350 1980.1200 3929.5050 1980.2000 ;
      RECT 0.0000 1979.7800 3929.5050 1980.1200 ;
      RECT 0.0000 1978.8400 3930.2400 1979.7800 ;
      RECT 0.0000 1978.4200 3929.5050 1978.8400 ;
      RECT 0.0000 1977.1400 3930.2400 1978.4200 ;
      RECT 0.0000 1976.8000 3929.5050 1977.1400 ;
      RECT 0.7350 1976.7200 3929.5050 1976.8000 ;
      RECT 0.7350 1976.3800 3930.2400 1976.7200 ;
      RECT 0.0000 1975.4400 3930.2400 1976.3800 ;
      RECT 0.0000 1975.0200 3929.5050 1975.4400 ;
      RECT 0.0000 1974.0800 3930.2400 1975.0200 ;
      RECT 0.0000 1973.6600 3929.5050 1974.0800 ;
      RECT 0.0000 1972.3800 3930.2400 1973.6600 ;
      RECT 0.0000 1971.9600 3929.5050 1972.3800 ;
      RECT 0.0000 1970.6800 3930.2400 1971.9600 ;
      RECT 0.0000 1970.2600 3929.5050 1970.6800 ;
      RECT 0.0000 1969.3200 3930.2400 1970.2600 ;
      RECT 0.0000 1968.9000 3929.5050 1969.3200 ;
      RECT 0.0000 1967.6200 3930.2400 1968.9000 ;
      RECT 0.0000 1967.2000 3929.5050 1967.6200 ;
      RECT 0.0000 1966.2600 3930.2400 1967.2000 ;
      RECT 0.0000 1965.8400 3929.5050 1966.2600 ;
      RECT 0.0000 1791.8400 3930.2400 1965.8400 ;
      RECT 0.7350 1791.4200 3930.2400 1791.8400 ;
      RECT 0.0000 1746.6200 3930.2400 1791.4200 ;
      RECT 0.7350 1746.2000 3929.5050 1746.6200 ;
      RECT 0.0000 1744.5800 3930.2400 1746.2000 ;
      RECT 0.0000 1744.1600 3929.5050 1744.5800 ;
      RECT 0.0000 1743.2200 3930.2400 1744.1600 ;
      RECT 0.0000 1742.8000 3929.5050 1743.2200 ;
      RECT 0.0000 1742.5400 3930.2400 1742.8000 ;
      RECT 0.7350 1742.1200 3930.2400 1742.5400 ;
      RECT 0.0000 1741.5200 3930.2400 1742.1200 ;
      RECT 0.0000 1741.1000 3929.5050 1741.5200 ;
      RECT 0.0000 1740.1600 3930.2400 1741.1000 ;
      RECT 0.0000 1739.7400 3929.5050 1740.1600 ;
      RECT 0.0000 1738.4600 3930.2400 1739.7400 ;
      RECT 0.7350 1738.0400 3929.5050 1738.4600 ;
      RECT 0.0000 1737.1000 3930.2400 1738.0400 ;
      RECT 0.0000 1736.6800 3929.5050 1737.1000 ;
      RECT 0.0000 1735.4000 3930.2400 1736.6800 ;
      RECT 0.0000 1735.0600 3929.5050 1735.4000 ;
      RECT 0.7350 1734.9800 3929.5050 1735.0600 ;
      RECT 0.7350 1734.6400 3930.2400 1734.9800 ;
      RECT 0.0000 1733.7000 3930.2400 1734.6400 ;
      RECT 0.0000 1733.2800 3929.5050 1733.7000 ;
      RECT 0.0000 1732.3400 3930.2400 1733.2800 ;
      RECT 0.0000 1731.9200 3929.5050 1732.3400 ;
      RECT 0.0000 1730.6400 3930.2400 1731.9200 ;
      RECT 0.7350 1730.2200 3929.5050 1730.6400 ;
      RECT 0.0000 1729.2800 3930.2400 1730.2200 ;
      RECT 0.0000 1728.8600 3929.5050 1729.2800 ;
      RECT 0.0000 1727.5800 3930.2400 1728.8600 ;
      RECT 0.0000 1727.1600 3929.5050 1727.5800 ;
      RECT 0.0000 1726.9000 3930.2400 1727.1600 ;
      RECT 0.7350 1726.4800 3930.2400 1726.9000 ;
      RECT 0.0000 1725.8800 3930.2400 1726.4800 ;
      RECT 0.0000 1725.4600 3929.5050 1725.8800 ;
      RECT 0.0000 1724.5200 3930.2400 1725.4600 ;
      RECT 0.0000 1724.1000 3929.5050 1724.5200 ;
      RECT 0.0000 1722.8200 3930.2400 1724.1000 ;
      RECT 0.0000 1722.4000 3929.5050 1722.8200 ;
      RECT 0.0000 1720.7800 3930.2400 1722.4000 ;
      RECT 0.0000 1720.3600 3929.5050 1720.7800 ;
      RECT 0.0000 1719.7600 3930.2400 1720.3600 ;
      RECT 0.0000 1719.3400 3929.5050 1719.7600 ;
      RECT 0.0000 1717.7200 3930.2400 1719.3400 ;
      RECT 0.0000 1717.3000 3929.5050 1717.7200 ;
      RECT 0.0000 1716.7000 3930.2400 1717.3000 ;
      RECT 0.0000 1716.2800 3929.5050 1716.7000 ;
      RECT 0.0000 1577.9800 3930.2400 1716.2800 ;
      RECT 0.7350 1577.5600 3930.2400 1577.9800 ;
      RECT 0.0000 1497.0600 3930.2400 1577.5600 ;
      RECT 0.7350 1496.7200 3930.2400 1497.0600 ;
      RECT 0.7350 1496.6400 3929.5050 1496.7200 ;
      RECT 0.0000 1496.3000 3929.5050 1496.6400 ;
      RECT 0.0000 1495.0200 3930.2400 1496.3000 ;
      RECT 0.0000 1494.6000 3929.5050 1495.0200 ;
      RECT 0.0000 1493.3200 3930.2400 1494.6000 ;
      RECT 0.0000 1492.9000 3929.5050 1493.3200 ;
      RECT 0.0000 1492.6400 3930.2400 1492.9000 ;
      RECT 0.7350 1492.2200 3930.2400 1492.6400 ;
      RECT 0.0000 1491.9600 3930.2400 1492.2200 ;
      RECT 0.0000 1491.5400 3929.5050 1491.9600 ;
      RECT 0.0000 1490.2600 3930.2400 1491.5400 ;
      RECT 0.0000 1489.8400 3929.5050 1490.2600 ;
      RECT 0.0000 1488.9000 3930.2400 1489.8400 ;
      RECT 0.7350 1488.5600 3930.2400 1488.9000 ;
      RECT 0.7350 1488.4800 3929.5050 1488.5600 ;
      RECT 0.0000 1488.1400 3929.5050 1488.4800 ;
      RECT 0.0000 1487.2000 3930.2400 1488.1400 ;
      RECT 0.0000 1486.7800 3929.5050 1487.2000 ;
      RECT 0.0000 1485.5000 3930.2400 1486.7800 ;
      RECT 0.0000 1485.1600 3929.5050 1485.5000 ;
      RECT 0.7350 1485.0800 3929.5050 1485.1600 ;
      RECT 0.7350 1484.7400 3930.2400 1485.0800 ;
      RECT 0.0000 1483.8000 3930.2400 1484.7400 ;
      RECT 0.0000 1483.3800 3929.5050 1483.8000 ;
      RECT 0.0000 1482.4400 3930.2400 1483.3800 ;
      RECT 0.0000 1482.0200 3929.5050 1482.4400 ;
      RECT 0.0000 1481.0800 3930.2400 1482.0200 ;
      RECT 0.7350 1480.7400 3930.2400 1481.0800 ;
      RECT 0.7350 1480.6600 3929.5050 1480.7400 ;
      RECT 0.0000 1480.3200 3929.5050 1480.6600 ;
      RECT 0.0000 1479.3800 3930.2400 1480.3200 ;
      RECT 0.0000 1478.9600 3929.5050 1479.3800 ;
      RECT 0.0000 1477.6800 3930.2400 1478.9600 ;
      RECT 0.0000 1477.3400 3929.5050 1477.6800 ;
      RECT 0.7350 1477.2600 3929.5050 1477.3400 ;
      RECT 0.7350 1476.9200 3930.2400 1477.2600 ;
      RECT 0.0000 1475.9800 3930.2400 1476.9200 ;
      RECT 0.0000 1475.5600 3929.5050 1475.9800 ;
      RECT 0.0000 1474.6200 3930.2400 1475.5600 ;
      RECT 0.0000 1474.2000 3929.5050 1474.6200 ;
      RECT 0.0000 1472.9200 3930.2400 1474.2000 ;
      RECT 0.0000 1472.5000 3929.5050 1472.9200 ;
      RECT 0.0000 1471.2200 3930.2400 1472.5000 ;
      RECT 0.0000 1470.8000 3929.5050 1471.2200 ;
      RECT 0.0000 1469.8600 3930.2400 1470.8000 ;
      RECT 0.0000 1469.4400 3929.5050 1469.8600 ;
      RECT 0.0000 1468.1600 3930.2400 1469.4400 ;
      RECT 0.0000 1467.7400 3929.5050 1468.1600 ;
      RECT 0.0000 1466.8000 3930.2400 1467.7400 ;
      RECT 0.0000 1466.3800 3929.5050 1466.8000 ;
      RECT 0.0000 1425.6600 3930.2400 1466.3800 ;
      RECT 0.7350 1425.2400 3930.2400 1425.6600 ;
      RECT 0.0000 1422.6000 3930.2400 1425.2400 ;
      RECT 0.7350 1422.1800 3930.2400 1422.6000 ;
      RECT 0.0000 1420.2200 3930.2400 1422.1800 ;
      RECT 0.7350 1419.8000 3930.2400 1420.2200 ;
      RECT 0.0000 1417.1600 3930.2400 1419.8000 ;
      RECT 0.7350 1416.7400 3930.2400 1417.1600 ;
      RECT 0.0000 1414.7800 3930.2400 1416.7400 ;
      RECT 0.7350 1414.3600 3930.2400 1414.7800 ;
      RECT 0.0000 1411.7200 3930.2400 1414.3600 ;
      RECT 0.7350 1411.3000 3930.2400 1411.7200 ;
      RECT 0.0000 1409.3400 3930.2400 1411.3000 ;
      RECT 0.7350 1408.9200 3930.2400 1409.3400 ;
      RECT 0.0000 1406.2800 3930.2400 1408.9200 ;
      RECT 0.7350 1405.8600 3930.2400 1406.2800 ;
      RECT 0.0000 1403.9000 3930.2400 1405.8600 ;
      RECT 0.7350 1403.4800 3930.2400 1403.9000 ;
      RECT 0.0000 1401.5200 3930.2400 1403.4800 ;
      RECT 0.7350 1401.1000 3930.2400 1401.5200 ;
      RECT 0.0000 1400.8400 3930.2400 1401.1000 ;
      RECT 0.7350 1400.4200 3930.2400 1400.8400 ;
      RECT 0.0000 1400.1600 3930.2400 1400.4200 ;
      RECT 0.7350 1399.7400 3930.2400 1400.1600 ;
      RECT 0.0000 1398.4600 3930.2400 1399.7400 ;
      RECT 0.7350 1398.0400 3930.2400 1398.4600 ;
      RECT 0.0000 1395.4000 3930.2400 1398.0400 ;
      RECT 0.7350 1394.9800 3930.2400 1395.4000 ;
      RECT 0.0000 1393.0200 3930.2400 1394.9800 ;
      RECT 0.7350 1392.6000 3930.2400 1393.0200 ;
      RECT 0.0000 1389.9600 3930.2400 1392.6000 ;
      RECT 0.7350 1389.5400 3930.2400 1389.9600 ;
      RECT 0.0000 1387.5800 3930.2400 1389.5400 ;
      RECT 0.7350 1387.1600 3930.2400 1387.5800 ;
      RECT 0.0000 1384.5200 3930.2400 1387.1600 ;
      RECT 0.7350 1384.1000 3930.2400 1384.5200 ;
      RECT 0.0000 1383.8400 3930.2400 1384.1000 ;
      RECT 0.7350 1383.4200 3930.2400 1383.8400 ;
      RECT 0.0000 1382.1400 3930.2400 1383.4200 ;
      RECT 0.7350 1381.7200 3930.2400 1382.1400 ;
      RECT 0.0000 1381.4600 3930.2400 1381.7200 ;
      RECT 0.7350 1381.0400 3930.2400 1381.4600 ;
      RECT 0.0000 1378.7400 3930.2400 1381.0400 ;
      RECT 0.7350 1378.3200 3930.2400 1378.7400 ;
      RECT 0.0000 1376.7000 3930.2400 1378.3200 ;
      RECT 0.7350 1376.2800 3930.2400 1376.7000 ;
      RECT 0.0000 1373.6400 3930.2400 1376.2800 ;
      RECT 0.7350 1373.2200 3930.2400 1373.6400 ;
      RECT 0.0000 1371.2600 3930.2400 1373.2200 ;
      RECT 0.7350 1370.8400 3930.2400 1371.2600 ;
      RECT 0.0000 1368.2000 3930.2400 1370.8400 ;
      RECT 0.7350 1367.7800 3930.2400 1368.2000 ;
      RECT 0.0000 1330.1200 3930.2400 1367.7800 ;
      RECT 0.7350 1329.7000 3930.2400 1330.1200 ;
      RECT 0.0000 1324.6800 3930.2400 1329.7000 ;
      RECT 0.7350 1324.2600 3930.2400 1324.6800 ;
      RECT 0.0000 1247.1600 3930.2400 1324.2600 ;
      RECT 0.7350 1246.8200 3930.2400 1247.1600 ;
      RECT 0.7350 1246.7400 3929.5050 1246.8200 ;
      RECT 0.0000 1246.4000 3929.5050 1246.7400 ;
      RECT 0.0000 1245.1200 3930.2400 1246.4000 ;
      RECT 0.0000 1244.7000 3929.5050 1245.1200 ;
      RECT 0.0000 1243.4200 3930.2400 1244.7000 ;
      RECT 0.0000 1243.0800 3929.5050 1243.4200 ;
      RECT 0.7350 1243.0000 3929.5050 1243.0800 ;
      RECT 0.7350 1242.6600 3930.2400 1243.0000 ;
      RECT 0.0000 1242.0600 3930.2400 1242.6600 ;
      RECT 0.0000 1241.6400 3929.5050 1242.0600 ;
      RECT 0.0000 1240.3600 3930.2400 1241.6400 ;
      RECT 0.0000 1239.9400 3929.5050 1240.3600 ;
      RECT 0.0000 1239.0000 3930.2400 1239.9400 ;
      RECT 0.7350 1238.6600 3930.2400 1239.0000 ;
      RECT 0.7350 1238.5800 3929.5050 1238.6600 ;
      RECT 0.0000 1238.2400 3929.5050 1238.5800 ;
      RECT 0.0000 1237.3000 3930.2400 1238.2400 ;
      RECT 0.0000 1236.8800 3929.5050 1237.3000 ;
      RECT 0.0000 1235.6000 3930.2400 1236.8800 ;
      RECT 0.0000 1235.2600 3929.5050 1235.6000 ;
      RECT 0.7350 1235.1800 3929.5050 1235.2600 ;
      RECT 0.7350 1234.8400 3930.2400 1235.1800 ;
      RECT 0.0000 1233.9000 3930.2400 1234.8400 ;
      RECT 0.0000 1233.4800 3929.5050 1233.9000 ;
      RECT 0.0000 1232.5400 3930.2400 1233.4800 ;
      RECT 0.0000 1232.1200 3929.5050 1232.5400 ;
      RECT 0.0000 1231.1800 3930.2400 1232.1200 ;
      RECT 0.7350 1230.8400 3930.2400 1231.1800 ;
      RECT 0.7350 1230.7600 3929.5050 1230.8400 ;
      RECT 0.0000 1230.4200 3929.5050 1230.7600 ;
      RECT 0.0000 1229.4800 3930.2400 1230.4200 ;
      RECT 0.0000 1229.0600 3929.5050 1229.4800 ;
      RECT 0.0000 1227.7800 3930.2400 1229.0600 ;
      RECT 0.0000 1227.4400 3929.5050 1227.7800 ;
      RECT 0.7350 1227.3600 3929.5050 1227.4400 ;
      RECT 0.7350 1227.0200 3930.2400 1227.3600 ;
      RECT 0.0000 1226.0800 3930.2400 1227.0200 ;
      RECT 0.0000 1225.6600 3929.5050 1226.0800 ;
      RECT 0.0000 1224.7200 3930.2400 1225.6600 ;
      RECT 0.0000 1224.3000 3929.5050 1224.7200 ;
      RECT 0.0000 1223.0200 3930.2400 1224.3000 ;
      RECT 0.0000 1222.6000 3929.5050 1223.0200 ;
      RECT 0.0000 1221.3200 3930.2400 1222.6000 ;
      RECT 0.0000 1220.9000 3929.5050 1221.3200 ;
      RECT 0.0000 1219.9600 3930.2400 1220.9000 ;
      RECT 0.0000 1219.5400 3929.5050 1219.9600 ;
      RECT 0.0000 1218.2600 3930.2400 1219.5400 ;
      RECT 0.0000 1217.8400 3929.5050 1218.2600 ;
      RECT 0.0000 1216.9000 3930.2400 1217.8400 ;
      RECT 0.0000 1216.4800 3929.5050 1216.9000 ;
      RECT 0.0000 997.2600 3930.2400 1216.4800 ;
      RECT 0.7350 996.9200 3930.2400 997.2600 ;
      RECT 0.7350 996.8400 3929.5050 996.9200 ;
      RECT 0.0000 996.5000 3929.5050 996.8400 ;
      RECT 0.0000 995.2200 3930.2400 996.5000 ;
      RECT 0.0000 994.8000 3929.5050 995.2200 ;
      RECT 0.0000 993.5200 3930.2400 994.8000 ;
      RECT 0.0000 993.1800 3929.5050 993.5200 ;
      RECT 0.7350 993.1000 3929.5050 993.1800 ;
      RECT 0.7350 992.7600 3930.2400 993.1000 ;
      RECT 0.0000 992.1600 3930.2400 992.7600 ;
      RECT 0.0000 991.7400 3929.5050 992.1600 ;
      RECT 0.0000 990.4600 3930.2400 991.7400 ;
      RECT 0.0000 990.0400 3929.5050 990.4600 ;
      RECT 0.0000 989.1000 3930.2400 990.0400 ;
      RECT 0.7350 988.7600 3930.2400 989.1000 ;
      RECT 0.7350 988.6800 3929.5050 988.7600 ;
      RECT 0.0000 988.3400 3929.5050 988.6800 ;
      RECT 0.0000 987.4000 3930.2400 988.3400 ;
      RECT 0.0000 986.9800 3929.5050 987.4000 ;
      RECT 0.0000 985.7000 3930.2400 986.9800 ;
      RECT 0.0000 985.3600 3929.5050 985.7000 ;
      RECT 0.7350 985.2800 3929.5050 985.3600 ;
      RECT 0.7350 984.9400 3930.2400 985.2800 ;
      RECT 0.0000 984.0000 3930.2400 984.9400 ;
      RECT 0.0000 983.5800 3929.5050 984.0000 ;
      RECT 0.0000 982.6400 3930.2400 983.5800 ;
      RECT 0.0000 982.2200 3929.5050 982.6400 ;
      RECT 0.0000 981.2800 3930.2400 982.2200 ;
      RECT 0.7350 980.9400 3930.2400 981.2800 ;
      RECT 0.7350 980.8600 3929.5050 980.9400 ;
      RECT 0.0000 980.5200 3929.5050 980.8600 ;
      RECT 0.0000 979.5800 3930.2400 980.5200 ;
      RECT 0.0000 979.1600 3929.5050 979.5800 ;
      RECT 0.0000 977.8800 3930.2400 979.1600 ;
      RECT 0.0000 977.5400 3929.5050 977.8800 ;
      RECT 0.7350 977.4600 3929.5050 977.5400 ;
      RECT 0.7350 977.1200 3930.2400 977.4600 ;
      RECT 0.0000 976.1800 3930.2400 977.1200 ;
      RECT 0.0000 975.7600 3929.5050 976.1800 ;
      RECT 0.0000 974.8200 3930.2400 975.7600 ;
      RECT 0.0000 974.4000 3929.5050 974.8200 ;
      RECT 0.0000 973.1200 3930.2400 974.4000 ;
      RECT 0.0000 972.7000 3929.5050 973.1200 ;
      RECT 0.0000 971.4200 3930.2400 972.7000 ;
      RECT 0.0000 971.0000 3929.5050 971.4200 ;
      RECT 0.0000 970.0600 3930.2400 971.0000 ;
      RECT 0.0000 969.6400 3929.5050 970.0600 ;
      RECT 0.0000 968.3600 3930.2400 969.6400 ;
      RECT 0.0000 967.9400 3929.5050 968.3600 ;
      RECT 0.0000 967.0000 3930.2400 967.9400 ;
      RECT 0.0000 966.5800 3929.5050 967.0000 ;
      RECT 0.0000 747.3600 3930.2400 966.5800 ;
      RECT 0.7350 747.0200 3930.2400 747.3600 ;
      RECT 0.7350 746.9400 3929.5050 747.0200 ;
      RECT 0.0000 746.6000 3929.5050 746.9400 ;
      RECT 0.0000 745.6600 3930.2400 746.6000 ;
      RECT 0.0000 745.2400 3929.5050 745.6600 ;
      RECT 0.0000 743.6200 3930.2400 745.2400 ;
      RECT 0.0000 743.2800 3929.5050 743.6200 ;
      RECT 0.7350 743.2000 3929.5050 743.2800 ;
      RECT 0.7350 742.8600 3930.2400 743.2000 ;
      RECT 0.0000 742.2600 3930.2400 742.8600 ;
      RECT 0.0000 741.8400 3929.5050 742.2600 ;
      RECT 0.0000 740.5600 3930.2400 741.8400 ;
      RECT 0.0000 740.1400 3929.5050 740.5600 ;
      RECT 0.0000 739.2000 3930.2400 740.1400 ;
      RECT 0.7350 738.8600 3930.2400 739.2000 ;
      RECT 0.7350 738.7800 3929.5050 738.8600 ;
      RECT 0.0000 738.4400 3929.5050 738.7800 ;
      RECT 0.0000 737.5000 3930.2400 738.4400 ;
      RECT 0.0000 737.0800 3929.5050 737.5000 ;
      RECT 0.0000 735.8000 3930.2400 737.0800 ;
      RECT 0.0000 735.4600 3929.5050 735.8000 ;
      RECT 0.7350 735.3800 3929.5050 735.4600 ;
      RECT 0.7350 735.0400 3930.2400 735.3800 ;
      RECT 0.0000 734.1000 3930.2400 735.0400 ;
      RECT 0.0000 733.6800 3929.5050 734.1000 ;
      RECT 0.0000 732.7400 3930.2400 733.6800 ;
      RECT 0.0000 732.3200 3929.5050 732.7400 ;
      RECT 0.0000 731.3800 3930.2400 732.3200 ;
      RECT 0.7350 731.0400 3930.2400 731.3800 ;
      RECT 0.7350 730.9600 3929.5050 731.0400 ;
      RECT 0.0000 730.6200 3929.5050 730.9600 ;
      RECT 0.0000 729.6800 3930.2400 730.6200 ;
      RECT 0.0000 729.2600 3929.5050 729.6800 ;
      RECT 0.0000 727.9800 3930.2400 729.2600 ;
      RECT 0.0000 727.6400 3929.5050 727.9800 ;
      RECT 0.7350 727.5600 3929.5050 727.6400 ;
      RECT 0.7350 727.2200 3930.2400 727.5600 ;
      RECT 0.0000 726.2800 3930.2400 727.2200 ;
      RECT 0.0000 725.8600 3929.5050 726.2800 ;
      RECT 0.0000 724.9200 3930.2400 725.8600 ;
      RECT 0.0000 724.5000 3929.5050 724.9200 ;
      RECT 0.0000 723.2200 3930.2400 724.5000 ;
      RECT 0.0000 722.8000 3929.5050 723.2200 ;
      RECT 0.0000 721.5200 3930.2400 722.8000 ;
      RECT 0.0000 721.1000 3929.5050 721.5200 ;
      RECT 0.0000 720.1600 3930.2400 721.1000 ;
      RECT 0.0000 719.7400 3929.5050 720.1600 ;
      RECT 0.0000 718.4600 3930.2400 719.7400 ;
      RECT 0.0000 718.0400 3929.5050 718.4600 ;
      RECT 0.0000 717.1000 3930.2400 718.0400 ;
      RECT 0.0000 716.6800 3929.5050 717.1000 ;
      RECT 0.0000 497.4600 3930.2400 716.6800 ;
      RECT 0.7350 497.1200 3930.2400 497.4600 ;
      RECT 0.7350 497.0400 3929.5050 497.1200 ;
      RECT 0.0000 496.7000 3929.5050 497.0400 ;
      RECT 0.0000 495.4200 3930.2400 496.7000 ;
      RECT 0.0000 495.0000 3929.5050 495.4200 ;
      RECT 0.0000 493.7200 3930.2400 495.0000 ;
      RECT 0.0000 493.3800 3929.5050 493.7200 ;
      RECT 0.7350 493.3000 3929.5050 493.3800 ;
      RECT 0.7350 492.9600 3930.2400 493.3000 ;
      RECT 0.0000 492.3600 3930.2400 492.9600 ;
      RECT 0.0000 491.9400 3929.5050 492.3600 ;
      RECT 0.0000 490.6600 3930.2400 491.9400 ;
      RECT 0.0000 490.2400 3929.5050 490.6600 ;
      RECT 0.0000 489.3000 3930.2400 490.2400 ;
      RECT 0.7350 488.9600 3930.2400 489.3000 ;
      RECT 0.7350 488.8800 3929.5050 488.9600 ;
      RECT 0.0000 488.5400 3929.5050 488.8800 ;
      RECT 0.0000 487.6000 3930.2400 488.5400 ;
      RECT 0.0000 487.1800 3929.5050 487.6000 ;
      RECT 0.0000 485.9000 3930.2400 487.1800 ;
      RECT 0.0000 485.5600 3929.5050 485.9000 ;
      RECT 0.7350 485.4800 3929.5050 485.5600 ;
      RECT 0.7350 485.1400 3930.2400 485.4800 ;
      RECT 0.0000 484.5400 3930.2400 485.1400 ;
      RECT 0.0000 484.1200 3929.5050 484.5400 ;
      RECT 0.0000 482.8400 3930.2400 484.1200 ;
      RECT 0.0000 482.4200 3929.5050 482.8400 ;
      RECT 0.0000 481.4800 3930.2400 482.4200 ;
      RECT 0.7350 481.0600 3929.5050 481.4800 ;
      RECT 0.0000 479.7800 3930.2400 481.0600 ;
      RECT 0.0000 479.3600 3929.5050 479.7800 ;
      RECT 0.0000 478.4200 3930.2400 479.3600 ;
      RECT 0.0000 478.0000 3929.5050 478.4200 ;
      RECT 0.0000 477.7400 3930.2400 478.0000 ;
      RECT 0.7350 477.3200 3930.2400 477.7400 ;
      RECT 0.0000 476.3800 3930.2400 477.3200 ;
      RECT 0.0000 475.9600 3929.5050 476.3800 ;
      RECT 0.0000 475.3600 3930.2400 475.9600 ;
      RECT 0.0000 474.9400 3929.5050 475.3600 ;
      RECT 0.0000 473.3200 3930.2400 474.9400 ;
      RECT 0.0000 472.9000 3929.5050 473.3200 ;
      RECT 0.0000 471.6200 3930.2400 472.9000 ;
      RECT 0.0000 471.2000 3929.5050 471.6200 ;
      RECT 0.0000 470.2600 3930.2400 471.2000 ;
      RECT 0.0000 469.8400 3929.5050 470.2600 ;
      RECT 0.0000 468.5600 3930.2400 469.8400 ;
      RECT 0.0000 468.1400 3929.5050 468.5600 ;
      RECT 0.0000 467.2000 3930.2400 468.1400 ;
      RECT 0.0000 466.7800 3929.5050 467.2000 ;
      RECT 0.0000 247.9000 3930.2400 466.7800 ;
      RECT 0.7350 247.5600 3930.2400 247.9000 ;
      RECT 0.7350 247.4800 3929.5050 247.5600 ;
      RECT 0.0000 247.1400 3929.5050 247.4800 ;
      RECT 0.0000 245.8600 3930.2400 247.1400 ;
      RECT 0.0000 245.4400 3929.5050 245.8600 ;
      RECT 0.0000 244.1600 3930.2400 245.4400 ;
      RECT 0.0000 243.7400 3929.5050 244.1600 ;
      RECT 0.0000 243.4800 3930.2400 243.7400 ;
      RECT 0.7350 243.0600 3930.2400 243.4800 ;
      RECT 0.0000 242.8000 3930.2400 243.0600 ;
      RECT 0.0000 242.3800 3929.5050 242.8000 ;
      RECT 0.0000 241.1000 3930.2400 242.3800 ;
      RECT 0.0000 240.6800 3929.5050 241.1000 ;
      RECT 0.0000 239.4000 3930.2400 240.6800 ;
      RECT 0.7350 239.0600 3930.2400 239.4000 ;
      RECT 0.7350 238.9800 3929.5050 239.0600 ;
      RECT 0.0000 238.6400 3929.5050 238.9800 ;
      RECT 0.0000 238.0400 3930.2400 238.6400 ;
      RECT 0.0000 237.6200 3929.5050 238.0400 ;
      RECT 0.0000 236.0000 3930.2400 237.6200 ;
      RECT 0.0000 235.6600 3929.5050 236.0000 ;
      RECT 0.7350 235.5800 3929.5050 235.6600 ;
      RECT 0.7350 235.2400 3930.2400 235.5800 ;
      RECT 0.0000 234.6400 3930.2400 235.2400 ;
      RECT 0.0000 234.2200 3929.5050 234.6400 ;
      RECT 0.0000 233.2800 3930.2400 234.2200 ;
      RECT 0.0000 232.8600 3929.5050 233.2800 ;
      RECT 0.0000 231.5800 3930.2400 232.8600 ;
      RECT 0.7350 231.1600 3929.5050 231.5800 ;
      RECT 0.0000 230.2200 3930.2400 231.1600 ;
      RECT 0.0000 229.8000 3929.5050 230.2200 ;
      RECT 0.0000 228.5200 3930.2400 229.8000 ;
      RECT 0.0000 228.1000 3929.5050 228.5200 ;
      RECT 0.0000 227.8400 3930.2400 228.1000 ;
      RECT 0.7350 227.4200 3930.2400 227.8400 ;
      RECT 0.0000 226.8200 3930.2400 227.4200 ;
      RECT 0.0000 226.4000 3929.5050 226.8200 ;
      RECT 0.0000 225.4600 3930.2400 226.4000 ;
      RECT 0.0000 225.0400 3929.5050 225.4600 ;
      RECT 0.0000 223.7600 3930.2400 225.0400 ;
      RECT 0.0000 223.3400 3929.5050 223.7600 ;
      RECT 0.0000 222.0600 3930.2400 223.3400 ;
      RECT 0.0000 221.6400 3929.5050 222.0600 ;
      RECT 0.0000 220.7000 3930.2400 221.6400 ;
      RECT 0.0000 220.2800 3929.5050 220.7000 ;
      RECT 0.0000 219.0000 3930.2400 220.2800 ;
      RECT 0.0000 218.5800 3929.5050 219.0000 ;
      RECT 0.0000 217.6400 3930.2400 218.5800 ;
      RECT 0.0000 217.2200 3929.5050 217.6400 ;
      RECT 0.0000 0.0000 3930.2400 217.2200 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 3930.2400 3930.0600 ;
    LAYER met3 ;
      RECT 0.0000 1403.9400 3930.2400 3930.0600 ;
      RECT 1.1000 1403.0400 3930.2400 1403.9400 ;
      RECT 0.0000 1400.8900 3930.2400 1403.0400 ;
      RECT 1.1000 1399.9900 3930.2400 1400.8900 ;
      RECT 0.0000 1395.4000 3930.2400 1399.9900 ;
      RECT 1.1000 1394.5000 3930.2400 1395.4000 ;
      RECT 0.0000 1392.9600 3930.2400 1394.5000 ;
      RECT 1.1000 1392.0600 3930.2400 1392.9600 ;
      RECT 0.0000 1389.9100 3930.2400 1392.0600 ;
      RECT 1.1000 1389.0100 3930.2400 1389.9100 ;
      RECT 0.0000 1388.0800 3930.2400 1389.0100 ;
      RECT 1.1000 1387.1800 3930.2400 1388.0800 ;
      RECT 0.0000 1385.0300 3930.2400 1387.1800 ;
      RECT 1.1000 1384.1300 3930.2400 1385.0300 ;
      RECT 0.0000 1382.5900 3930.2400 1384.1300 ;
      RECT 1.1000 1381.6900 3930.2400 1382.5900 ;
      RECT 0.0000 1368.5600 3930.2400 1381.6900 ;
      RECT 1.1000 1367.6600 3930.2400 1368.5600 ;
      RECT 0.0000 0.0000 3930.2400 1367.6600 ;
    LAYER met4 ;
      RECT 0.0000 3928.4600 3930.2400 3930.0600 ;
      RECT 6.4000 3928.3600 3923.8400 3928.4600 ;
      RECT 3766.3800 3922.4600 3923.8400 3928.3600 ;
      RECT 6.4000 3922.4600 120.8800 3928.3600 ;
      RECT 3766.3800 3922.3600 3917.8400 3922.4600 ;
      RECT 3525.9200 3922.3600 3763.7800 3928.3600 ;
      RECT 3285.4600 3922.3600 3523.3200 3928.3600 ;
      RECT 3045.0000 3922.3600 3282.8600 3928.3600 ;
      RECT 2804.5400 3922.3600 3042.4000 3928.3600 ;
      RECT 2564.0800 3922.3600 2801.9400 3928.3600 ;
      RECT 2323.6200 3922.3600 2561.4800 3928.3600 ;
      RECT 2083.1600 3922.3600 2321.0200 3928.3600 ;
      RECT 1842.7000 3922.3600 2080.5600 3928.3600 ;
      RECT 1602.2400 3922.3600 1840.1000 3928.3600 ;
      RECT 1361.7800 3922.3600 1599.6400 3928.3600 ;
      RECT 1121.3200 3922.3600 1359.1800 3928.3600 ;
      RECT 880.8600 3922.3600 1118.7200 3928.3600 ;
      RECT 640.4000 3922.3600 878.2600 3928.3600 ;
      RECT 399.9400 3922.3600 637.8000 3928.3600 ;
      RECT 159.3800 3922.3600 397.3400 3928.3600 ;
      RECT 12.4000 3922.3600 120.8800 3922.4600 ;
      RECT 3529.9200 3913.2400 3763.7800 3922.3600 ;
      RECT 3525.9200 3913.2400 3527.3200 3922.3600 ;
      RECT 3289.4600 3913.2400 3523.3200 3922.3600 ;
      RECT 3285.4600 3913.2400 3286.8600 3922.3600 ;
      RECT 3049.0000 3913.2400 3282.8600 3922.3600 ;
      RECT 3045.0000 3913.2400 3046.4000 3922.3600 ;
      RECT 2808.5400 3913.2400 3042.4000 3922.3600 ;
      RECT 2804.5400 3913.2400 2805.9400 3922.3600 ;
      RECT 2568.0800 3913.2400 2801.9400 3922.3600 ;
      RECT 2564.0800 3913.2400 2565.4800 3922.3600 ;
      RECT 2327.6200 3913.2400 2561.4800 3922.3600 ;
      RECT 2323.6200 3913.2400 2325.0200 3922.3600 ;
      RECT 2087.1600 3913.2400 2321.0200 3922.3600 ;
      RECT 2083.1600 3913.2400 2084.5600 3922.3600 ;
      RECT 1846.7000 3913.2400 2080.5600 3922.3600 ;
      RECT 1842.7000 3913.2400 1844.1000 3922.3600 ;
      RECT 1606.2400 3913.2400 1840.1000 3922.3600 ;
      RECT 1602.2400 3913.2400 1603.6400 3922.3600 ;
      RECT 1365.7800 3913.2400 1599.6400 3922.3600 ;
      RECT 1361.7800 3913.2400 1363.1800 3922.3600 ;
      RECT 1125.3200 3913.2400 1359.1800 3922.3600 ;
      RECT 1121.3200 3913.2400 1122.7200 3922.3600 ;
      RECT 884.8600 3913.2400 1118.7200 3922.3600 ;
      RECT 880.8600 3913.2400 882.2600 3922.3600 ;
      RECT 644.4000 3913.2400 878.2600 3922.3600 ;
      RECT 640.4000 3913.2400 641.8000 3922.3600 ;
      RECT 403.9400 3913.2400 637.8000 3922.3600 ;
      RECT 399.9400 3913.2400 401.3400 3922.3600 ;
      RECT 163.3800 3913.2400 397.3400 3922.3600 ;
      RECT 159.3800 3913.2400 160.7800 3922.3600 ;
      RECT 3535.5800 3913.1400 3763.7800 3913.2400 ;
      RECT 3295.1200 3913.1400 3523.3200 3913.2400 ;
      RECT 3054.6600 3913.1400 3282.8600 3913.2400 ;
      RECT 2814.2000 3913.1400 3042.4000 3913.2400 ;
      RECT 2573.7400 3913.1400 2801.9400 3913.2400 ;
      RECT 2333.2800 3913.1400 2561.4800 3913.2400 ;
      RECT 2092.8200 3913.1400 2321.0200 3913.2400 ;
      RECT 1852.3600 3913.1400 2080.5600 3913.2400 ;
      RECT 1611.9000 3913.1400 1840.1000 3913.2400 ;
      RECT 1371.4400 3913.1400 1599.6400 3913.2400 ;
      RECT 1130.9800 3913.1400 1359.1800 3913.2400 ;
      RECT 890.5200 3913.1400 1118.7200 3913.2400 ;
      RECT 650.0600 3913.1400 878.2600 3913.2400 ;
      RECT 409.6000 3913.1400 637.8000 3913.2400 ;
      RECT 169.1400 3913.1400 397.3400 3913.2400 ;
      RECT 3536.4800 3910.5400 3763.7800 3913.1400 ;
      RECT 3296.0200 3910.5400 3523.3200 3913.1400 ;
      RECT 3055.5600 3910.5400 3282.8600 3913.1400 ;
      RECT 2815.1000 3910.5400 3042.4000 3913.1400 ;
      RECT 2574.6400 3910.5400 2801.9400 3913.1400 ;
      RECT 2334.1800 3910.5400 2561.4800 3913.1400 ;
      RECT 2093.7200 3910.5400 2321.0200 3913.1400 ;
      RECT 1853.2600 3910.5400 2080.5600 3913.1400 ;
      RECT 1612.8000 3910.5400 1840.1000 3913.1400 ;
      RECT 1372.3400 3910.5400 1599.6400 3913.1400 ;
      RECT 1131.8800 3910.5400 1359.1800 3913.1400 ;
      RECT 891.4200 3910.5400 1118.7200 3913.1400 ;
      RECT 650.9600 3910.5400 878.2600 3913.1400 ;
      RECT 410.5000 3910.5400 637.8000 3913.1400 ;
      RECT 170.0400 3910.5400 397.3400 3913.1400 ;
      RECT 3535.5800 3910.4400 3763.7800 3910.5400 ;
      RECT 3525.9200 3910.4400 3527.2200 3913.2400 ;
      RECT 3295.1200 3910.4400 3523.3200 3910.5400 ;
      RECT 3285.4600 3910.4400 3286.7600 3913.2400 ;
      RECT 3054.6600 3910.4400 3282.8600 3910.5400 ;
      RECT 3045.0000 3910.4400 3046.3000 3913.2400 ;
      RECT 2814.2000 3910.4400 3042.4000 3910.5400 ;
      RECT 2804.5400 3910.4400 2805.8400 3913.2400 ;
      RECT 2573.7400 3910.4400 2801.9400 3910.5400 ;
      RECT 2564.0800 3910.4400 2565.3800 3913.2400 ;
      RECT 2333.2800 3910.4400 2561.4800 3910.5400 ;
      RECT 2323.6200 3910.4400 2324.9200 3913.2400 ;
      RECT 2092.8200 3910.4400 2321.0200 3910.5400 ;
      RECT 2083.1600 3910.4400 2084.4600 3913.2400 ;
      RECT 1852.3600 3910.4400 2080.5600 3910.5400 ;
      RECT 1842.7000 3910.4400 1844.0000 3913.2400 ;
      RECT 1611.9000 3910.4400 1840.1000 3910.5400 ;
      RECT 1602.2400 3910.4400 1603.5400 3913.2400 ;
      RECT 1371.4400 3910.4400 1599.6400 3910.5400 ;
      RECT 1361.7800 3910.4400 1363.0800 3913.2400 ;
      RECT 1130.9800 3910.4400 1359.1800 3910.5400 ;
      RECT 1121.3200 3910.4400 1122.6200 3913.2400 ;
      RECT 890.5200 3910.4400 1118.7200 3910.5400 ;
      RECT 880.8600 3910.4400 882.1600 3913.2400 ;
      RECT 650.0600 3910.4400 878.2600 3910.5400 ;
      RECT 640.4000 3910.4400 641.7000 3913.2400 ;
      RECT 409.6000 3910.4400 637.8000 3910.5400 ;
      RECT 399.9400 3910.4400 401.2400 3913.2400 ;
      RECT 169.1400 3910.4400 397.3400 3910.5400 ;
      RECT 159.3800 3910.4400 160.6800 3913.2400 ;
      RECT 3529.9200 3891.2100 3763.7800 3910.4400 ;
      RECT 3289.4600 3891.2100 3523.3200 3910.4400 ;
      RECT 3049.0000 3891.2100 3282.8600 3910.4400 ;
      RECT 2808.5400 3891.2100 3042.4000 3910.4400 ;
      RECT 2568.0800 3891.2100 2801.9400 3910.4400 ;
      RECT 2327.6200 3891.2100 2561.4800 3910.4400 ;
      RECT 2087.1600 3891.2100 2321.0200 3910.4400 ;
      RECT 1846.7000 3891.2100 2080.5600 3910.4400 ;
      RECT 1606.2400 3891.2100 1840.1000 3910.4400 ;
      RECT 1365.7800 3891.2100 1599.6400 3910.4400 ;
      RECT 1125.3200 3891.2100 1359.1800 3910.4400 ;
      RECT 884.8600 3891.2100 1118.7200 3910.4400 ;
      RECT 644.4000 3891.2100 878.2600 3910.4400 ;
      RECT 403.9400 3891.2100 637.8000 3910.4400 ;
      RECT 163.3800 3891.2100 397.3400 3910.4400 ;
      RECT 3756.8200 3888.6100 3763.7800 3891.2100 ;
      RECT 3529.9200 3888.6100 3754.2200 3891.2100 ;
      RECT 3516.3600 3888.6100 3523.3200 3891.2100 ;
      RECT 3289.4600 3888.6100 3513.7600 3891.2100 ;
      RECT 3275.9000 3888.6100 3282.8600 3891.2100 ;
      RECT 3049.0000 3888.6100 3273.3000 3891.2100 ;
      RECT 3035.4400 3888.6100 3042.4000 3891.2100 ;
      RECT 2808.5400 3888.6100 3032.8400 3891.2100 ;
      RECT 2794.9800 3888.6100 2801.9400 3891.2100 ;
      RECT 2568.0800 3888.6100 2792.3800 3891.2100 ;
      RECT 2554.5200 3888.6100 2561.4800 3891.2100 ;
      RECT 2327.6200 3888.6100 2551.9200 3891.2100 ;
      RECT 2314.0600 3888.6100 2321.0200 3891.2100 ;
      RECT 2087.1600 3888.6100 2311.4600 3891.2100 ;
      RECT 2073.6000 3888.6100 2080.5600 3891.2100 ;
      RECT 1846.7000 3888.6100 2071.0000 3891.2100 ;
      RECT 1833.1400 3888.6100 1840.1000 3891.2100 ;
      RECT 1606.2400 3888.6100 1830.5400 3891.2100 ;
      RECT 1592.6800 3888.6100 1599.6400 3891.2100 ;
      RECT 1365.7800 3888.6100 1590.0800 3891.2100 ;
      RECT 1352.2200 3888.6100 1359.1800 3891.2100 ;
      RECT 1125.3200 3888.6100 1349.6200 3891.2100 ;
      RECT 1111.7600 3888.6100 1118.7200 3891.2100 ;
      RECT 884.8600 3888.6100 1109.1600 3891.2100 ;
      RECT 871.3000 3888.6100 878.2600 3891.2100 ;
      RECT 644.4000 3888.6100 868.7000 3891.2100 ;
      RECT 630.8400 3888.6100 637.8000 3891.2100 ;
      RECT 403.9400 3888.6100 628.2400 3891.2100 ;
      RECT 390.3800 3888.6100 397.3400 3891.2100 ;
      RECT 163.3800 3888.6100 387.7800 3891.2100 ;
      RECT 3770.3800 3867.1400 3917.8400 3922.3600 ;
      RECT 3529.9200 3643.7300 3763.7800 3888.6100 ;
      RECT 3289.4600 3643.7300 3523.3200 3888.6100 ;
      RECT 3049.0000 3643.7300 3282.8600 3888.6100 ;
      RECT 2808.5400 3643.7300 3042.4000 3888.6100 ;
      RECT 2327.6200 3643.7300 2561.4800 3888.6100 ;
      RECT 2087.1600 3643.7300 2321.0200 3888.6100 ;
      RECT 1846.7000 3643.7300 2080.5600 3888.6100 ;
      RECT 1606.2400 3643.7300 1840.1000 3888.6100 ;
      RECT 1365.7800 3643.7300 1599.6400 3888.6100 ;
      RECT 1125.3200 3643.7300 1359.1800 3888.6100 ;
      RECT 884.8600 3643.7300 1118.7200 3888.6100 ;
      RECT 644.4000 3643.7300 878.2600 3888.6100 ;
      RECT 403.9400 3643.7300 637.8000 3888.6100 ;
      RECT 163.3800 3643.7300 397.3400 3888.6100 ;
      RECT 159.3800 3642.5900 160.7800 3910.4400 ;
      RECT 123.4800 3642.5900 156.7800 3928.3600 ;
      RECT 123.4800 3642.4900 150.4400 3642.5900 ;
      RECT 3816.2800 3642.3300 3817.6800 3867.1400 ;
      RECT 3780.3800 3642.3300 3813.6800 3867.1400 ;
      RECT 3780.3800 3642.2300 3807.3400 3642.3300 ;
      RECT 123.4800 3640.3900 149.7900 3642.4900 ;
      RECT 159.4800 3640.2900 160.7800 3642.5900 ;
      RECT 123.4800 3640.2900 150.4400 3640.3900 ;
      RECT 3780.3800 3640.1300 3806.6900 3642.2300 ;
      RECT 3816.3800 3640.0300 3817.6800 3642.3300 ;
      RECT 3780.3800 3640.0300 3807.3400 3640.1300 ;
      RECT 123.4800 3639.9900 156.7800 3640.2900 ;
      RECT 3780.3800 3639.8300 3813.6800 3640.0300 ;
      RECT 3776.3800 3639.8300 3777.7800 3867.1400 ;
      RECT 3784.2200 3639.7300 3813.6800 3639.8300 ;
      RECT 3529.9200 3639.3300 3753.7200 3643.7300 ;
      RECT 3525.9200 3639.3300 3527.3200 3910.4400 ;
      RECT 3289.4600 3639.3300 3513.2600 3643.7300 ;
      RECT 3285.4600 3639.3300 3286.8600 3910.4400 ;
      RECT 3049.0000 3639.3300 3272.8000 3643.7300 ;
      RECT 3045.0000 3639.3300 3046.4000 3910.4400 ;
      RECT 2808.5400 3639.3300 3032.3400 3643.7300 ;
      RECT 2804.5400 3639.3300 2805.9400 3910.4400 ;
      RECT 2327.6200 3639.3300 2551.4200 3643.7300 ;
      RECT 2323.6200 3639.3300 2325.0200 3910.4400 ;
      RECT 2087.1600 3639.3300 2310.9600 3643.7300 ;
      RECT 2083.1600 3639.3300 2084.5600 3910.4400 ;
      RECT 1846.7000 3639.3300 2070.5000 3643.7300 ;
      RECT 1842.7000 3639.3300 1844.1000 3910.4400 ;
      RECT 1606.2400 3639.3300 1830.0400 3643.7300 ;
      RECT 1602.2400 3639.3300 1603.6400 3910.4400 ;
      RECT 1365.7800 3639.3300 1589.5800 3643.7300 ;
      RECT 1361.7800 3639.3300 1363.1800 3910.4400 ;
      RECT 1125.3200 3639.3300 1349.1200 3643.7300 ;
      RECT 1121.3200 3639.3300 1122.7200 3910.4400 ;
      RECT 884.8600 3639.3300 1108.6600 3643.7300 ;
      RECT 880.8600 3639.3300 882.2600 3910.4400 ;
      RECT 644.4000 3639.3300 868.2000 3643.7300 ;
      RECT 640.4000 3639.3300 641.8000 3910.4400 ;
      RECT 403.9400 3639.3300 627.7400 3643.7300 ;
      RECT 399.9400 3639.3300 401.3400 3910.4400 ;
      RECT 163.3800 3639.3300 387.2800 3643.7300 ;
      RECT 159.3800 3639.3300 160.7800 3640.2900 ;
      RECT 3535.0800 3639.2300 3753.7200 3639.3300 ;
      RECT 3294.6200 3639.2300 3513.2600 3639.3300 ;
      RECT 3054.1600 3639.2300 3272.8000 3639.3300 ;
      RECT 2813.7000 3639.2300 3032.3400 3639.3300 ;
      RECT 2332.7800 3639.2300 2551.4200 3639.3300 ;
      RECT 2092.3200 3639.2300 2310.9600 3639.3300 ;
      RECT 1851.8600 3639.2300 2070.5000 3639.3300 ;
      RECT 1611.4000 3639.2300 1830.0400 3639.3300 ;
      RECT 1370.9400 3639.2300 1589.5800 3639.3300 ;
      RECT 1130.4800 3639.2300 1349.1200 3639.3300 ;
      RECT 890.0200 3639.2300 1108.6600 3639.3300 ;
      RECT 649.5600 3639.2300 868.2000 3639.3300 ;
      RECT 409.1000 3639.2300 627.7400 3639.3300 ;
      RECT 168.6400 3639.2300 387.2800 3639.3300 ;
      RECT 156.3100 3637.8900 156.7800 3639.9900 ;
      RECT 123.4800 3637.8900 151.7050 3639.9900 ;
      RECT 3784.8700 3637.6300 3813.6800 3639.7300 ;
      RECT 3784.2200 3637.5300 3813.6800 3637.6300 ;
      RECT 3776.3800 3637.5300 3777.6800 3639.8300 ;
      RECT 3536.4800 3636.6300 3753.7200 3639.2300 ;
      RECT 3296.0200 3636.6300 3513.2600 3639.2300 ;
      RECT 3055.5600 3636.6300 3272.8000 3639.2300 ;
      RECT 2815.1000 3636.6300 3032.3400 3639.2300 ;
      RECT 2334.1800 3636.6300 2551.4200 3639.2300 ;
      RECT 2093.7200 3636.6300 2310.9600 3639.2300 ;
      RECT 1853.2600 3636.6300 2070.5000 3639.2300 ;
      RECT 1612.8000 3636.6300 1830.0400 3639.2300 ;
      RECT 1372.3400 3636.6300 1589.5800 3639.2300 ;
      RECT 1131.8800 3636.6300 1349.1200 3639.2300 ;
      RECT 891.4200 3636.6300 1108.6600 3639.2300 ;
      RECT 650.9600 3636.6300 868.2000 3639.2300 ;
      RECT 410.5000 3636.6300 627.7400 3639.2300 ;
      RECT 170.0400 3636.6300 387.2800 3639.2300 ;
      RECT 3535.0800 3636.5300 3753.7200 3636.6300 ;
      RECT 3525.9200 3636.5300 3527.2200 3639.3300 ;
      RECT 3294.6200 3636.5300 3513.2600 3636.6300 ;
      RECT 3285.4600 3636.5300 3286.7600 3639.3300 ;
      RECT 3054.1600 3636.5300 3272.8000 3636.6300 ;
      RECT 3045.0000 3636.5300 3046.3000 3639.3300 ;
      RECT 2813.7000 3636.5300 3032.3400 3636.6300 ;
      RECT 2804.5400 3636.5300 2805.8400 3639.3300 ;
      RECT 2332.7800 3636.5300 2551.4200 3636.6300 ;
      RECT 2323.6200 3636.5300 2324.9200 3639.3300 ;
      RECT 2092.3200 3636.5300 2310.9600 3636.6300 ;
      RECT 2083.1600 3636.5300 2084.4600 3639.3300 ;
      RECT 1851.8600 3636.5300 2070.5000 3636.6300 ;
      RECT 1842.7000 3636.5300 1844.0000 3639.3300 ;
      RECT 1611.4000 3636.5300 1830.0400 3636.6300 ;
      RECT 1602.2400 3636.5300 1603.5400 3639.3300 ;
      RECT 1370.9400 3636.5300 1589.5800 3636.6300 ;
      RECT 1361.7800 3636.5300 1363.0800 3639.3300 ;
      RECT 1130.4800 3636.5300 1349.1200 3636.6300 ;
      RECT 1121.3200 3636.5300 1122.6200 3639.3300 ;
      RECT 890.0200 3636.5300 1108.6600 3636.6300 ;
      RECT 880.8600 3636.5300 882.1600 3639.3300 ;
      RECT 649.5600 3636.5300 868.2000 3636.6300 ;
      RECT 640.4000 3636.5300 641.7000 3639.3300 ;
      RECT 409.1000 3636.5300 627.7400 3636.6300 ;
      RECT 399.9400 3636.5300 401.2400 3639.3300 ;
      RECT 168.6400 3636.5300 387.2800 3636.6300 ;
      RECT 159.3800 3636.5300 160.6800 3639.3300 ;
      RECT 3776.3800 3632.7000 3777.7800 3637.5300 ;
      RECT 3770.3800 3632.7000 3773.7800 3867.1400 ;
      RECT 3816.2800 3630.7000 3817.6800 3640.0300 ;
      RECT 3780.3800 3630.7000 3813.6800 3637.5300 ;
      RECT 3756.3200 3630.7000 3763.7800 3643.7300 ;
      RECT 3529.9200 3630.7000 3753.7200 3636.5300 ;
      RECT 3515.8600 3630.7000 3523.3200 3643.7300 ;
      RECT 3289.4600 3630.7000 3513.2600 3636.5300 ;
      RECT 3275.4000 3630.7000 3282.8600 3643.7300 ;
      RECT 3049.0000 3630.7000 3272.8000 3636.5300 ;
      RECT 3034.9400 3630.7000 3042.4000 3643.7300 ;
      RECT 2808.5400 3630.7000 3032.3400 3636.5300 ;
      RECT 2554.0200 3630.7000 2561.4800 3643.7300 ;
      RECT 2327.6200 3630.7000 2551.4200 3636.5300 ;
      RECT 2313.5600 3630.7000 2321.0200 3643.7300 ;
      RECT 2087.1600 3630.7000 2310.9600 3636.5300 ;
      RECT 2073.1000 3630.7000 2080.5600 3643.7300 ;
      RECT 1846.7000 3630.7000 2070.5000 3636.5300 ;
      RECT 1832.6400 3630.7000 1840.1000 3643.7300 ;
      RECT 1606.2400 3630.7000 1830.0400 3636.5300 ;
      RECT 1592.1800 3630.7000 1599.6400 3643.7300 ;
      RECT 1365.7800 3630.7000 1589.5800 3636.5300 ;
      RECT 1351.7200 3630.7000 1359.1800 3643.7300 ;
      RECT 1125.3200 3630.7000 1349.1200 3636.5300 ;
      RECT 1111.2600 3630.7000 1118.7200 3643.7300 ;
      RECT 884.8600 3630.7000 1108.6600 3636.5300 ;
      RECT 870.8000 3630.7000 878.2600 3643.7300 ;
      RECT 644.4000 3630.7000 868.2000 3636.5300 ;
      RECT 630.3400 3630.7000 637.8000 3643.7300 ;
      RECT 403.9400 3630.7000 627.7400 3636.5300 ;
      RECT 389.8800 3630.7000 397.3400 3643.7300 ;
      RECT 163.3800 3630.7000 387.2800 3636.5300 ;
      RECT 3820.2800 3626.7000 3917.8400 3867.1400 ;
      RECT 3780.3800 3626.7000 3817.6800 3630.7000 ;
      RECT 3770.3800 3626.7000 3777.7800 3632.7000 ;
      RECT 3770.3800 3617.3000 3917.8400 3626.7000 ;
      RECT 3529.9200 3393.8900 3763.7800 3630.7000 ;
      RECT 3289.4600 3393.8900 3523.3200 3630.7000 ;
      RECT 3049.0000 3393.8900 3282.8600 3630.7000 ;
      RECT 2808.5400 3393.8900 3042.4000 3630.7000 ;
      RECT 2568.0800 3393.8900 2801.9400 3888.6100 ;
      RECT 2327.6200 3393.8900 2561.4800 3630.7000 ;
      RECT 2087.1600 3393.8900 2321.0200 3630.7000 ;
      RECT 1846.7000 3393.8900 2080.5600 3630.7000 ;
      RECT 1606.2400 3393.8900 1840.1000 3630.7000 ;
      RECT 1365.7800 3393.8900 1599.6400 3630.7000 ;
      RECT 1125.3200 3393.8900 1359.1800 3630.7000 ;
      RECT 884.8600 3393.8900 1118.7200 3630.7000 ;
      RECT 644.4000 3393.8900 878.2600 3630.7000 ;
      RECT 403.9400 3393.8900 637.8000 3630.7000 ;
      RECT 163.3800 3393.8900 397.3400 3630.7000 ;
      RECT 159.3800 3392.7500 160.7800 3636.5300 ;
      RECT 123.4800 3392.7500 156.7800 3637.8900 ;
      RECT 123.4800 3392.6500 150.4400 3392.7500 ;
      RECT 3816.2800 3392.4900 3817.6800 3617.3000 ;
      RECT 3780.3800 3392.4900 3813.6800 3617.3000 ;
      RECT 3780.3800 3392.3900 3807.3400 3392.4900 ;
      RECT 123.4800 3390.5500 149.7900 3392.6500 ;
      RECT 159.4800 3390.4500 160.7800 3392.7500 ;
      RECT 123.4800 3390.4500 150.4400 3390.5500 ;
      RECT 3780.3800 3390.2900 3806.6900 3392.3900 ;
      RECT 3816.3800 3390.1900 3817.6800 3392.4900 ;
      RECT 3780.3800 3390.1900 3807.3400 3390.2900 ;
      RECT 123.4800 3390.1500 156.7800 3390.4500 ;
      RECT 3780.3800 3389.9900 3813.6800 3390.1900 ;
      RECT 3776.3800 3389.9900 3777.7800 3617.3000 ;
      RECT 3784.2200 3389.8900 3813.6800 3389.9900 ;
      RECT 3529.9200 3389.4900 3753.7200 3393.8900 ;
      RECT 3525.9200 3389.4900 3527.3200 3636.5300 ;
      RECT 3289.4600 3389.4900 3513.2600 3393.8900 ;
      RECT 3285.4600 3389.4900 3286.8600 3636.5300 ;
      RECT 3049.0000 3389.4900 3272.8000 3393.8900 ;
      RECT 3045.0000 3389.4900 3046.4000 3636.5300 ;
      RECT 2808.5400 3389.4900 3032.3400 3393.8900 ;
      RECT 2804.5400 3389.4900 2805.9400 3636.5300 ;
      RECT 2568.0800 3389.4900 2791.8800 3393.8900 ;
      RECT 2564.0800 3389.4900 2565.4800 3910.4400 ;
      RECT 2327.6200 3389.4900 2551.4200 3393.8900 ;
      RECT 2323.6200 3389.4900 2325.0200 3636.5300 ;
      RECT 2087.1600 3389.4900 2310.9600 3393.8900 ;
      RECT 2083.1600 3389.4900 2084.5600 3636.5300 ;
      RECT 1846.7000 3389.4900 2070.5000 3393.8900 ;
      RECT 1842.7000 3389.4900 1844.1000 3636.5300 ;
      RECT 1606.2400 3389.4900 1830.0400 3393.8900 ;
      RECT 1602.2400 3389.4900 1603.6400 3636.5300 ;
      RECT 1365.7800 3389.4900 1589.5800 3393.8900 ;
      RECT 1361.7800 3389.4900 1363.1800 3636.5300 ;
      RECT 1125.3200 3389.4900 1349.1200 3393.8900 ;
      RECT 1121.3200 3389.4900 1122.7200 3636.5300 ;
      RECT 884.8600 3389.4900 1108.6600 3393.8900 ;
      RECT 880.8600 3389.4900 882.2600 3636.5300 ;
      RECT 644.4000 3389.4900 868.2000 3393.8900 ;
      RECT 640.4000 3389.4900 641.8000 3636.5300 ;
      RECT 403.9400 3389.4900 627.7400 3393.8900 ;
      RECT 399.9400 3389.4900 401.3400 3636.5300 ;
      RECT 163.3800 3389.4900 387.2800 3393.8900 ;
      RECT 159.3800 3389.4900 160.7800 3390.4500 ;
      RECT 3535.0800 3389.3900 3753.7200 3389.4900 ;
      RECT 3294.6200 3389.3900 3513.2600 3389.4900 ;
      RECT 3054.1600 3389.3900 3272.8000 3389.4900 ;
      RECT 2813.7000 3389.3900 3032.3400 3389.4900 ;
      RECT 2573.2400 3389.3900 2791.8800 3389.4900 ;
      RECT 2332.7800 3389.3900 2551.4200 3389.4900 ;
      RECT 2092.3200 3389.3900 2310.9600 3389.4900 ;
      RECT 1851.8600 3389.3900 2070.5000 3389.4900 ;
      RECT 1611.4000 3389.3900 1830.0400 3389.4900 ;
      RECT 1370.9400 3389.3900 1589.5800 3389.4900 ;
      RECT 1130.4800 3389.3900 1349.1200 3389.4900 ;
      RECT 890.0200 3389.3900 1108.6600 3389.4900 ;
      RECT 649.5600 3389.3900 868.2000 3389.4900 ;
      RECT 409.1000 3389.3900 627.7400 3389.4900 ;
      RECT 168.6400 3389.3900 387.2800 3389.4900 ;
      RECT 156.3100 3388.0500 156.7800 3390.1500 ;
      RECT 123.4800 3388.0500 151.7050 3390.1500 ;
      RECT 3784.8700 3387.7900 3813.6800 3389.8900 ;
      RECT 3784.2200 3387.6900 3813.6800 3387.7900 ;
      RECT 3776.3800 3387.6900 3777.6800 3389.9900 ;
      RECT 3536.4800 3386.7900 3753.7200 3389.3900 ;
      RECT 3296.0200 3386.7900 3513.2600 3389.3900 ;
      RECT 3055.5600 3386.7900 3272.8000 3389.3900 ;
      RECT 2815.1000 3386.7900 3032.3400 3389.3900 ;
      RECT 2574.6400 3386.7900 2791.8800 3389.3900 ;
      RECT 2334.1800 3386.7900 2551.4200 3389.3900 ;
      RECT 2093.7200 3386.7900 2310.9600 3389.3900 ;
      RECT 1853.2600 3386.7900 2070.5000 3389.3900 ;
      RECT 1612.8000 3386.7900 1830.0400 3389.3900 ;
      RECT 1372.3400 3386.7900 1589.5800 3389.3900 ;
      RECT 1131.8800 3386.7900 1349.1200 3389.3900 ;
      RECT 891.4200 3386.7900 1108.6600 3389.3900 ;
      RECT 650.9600 3386.7900 868.2000 3389.3900 ;
      RECT 410.5000 3386.7900 627.7400 3389.3900 ;
      RECT 170.0400 3386.7900 387.2800 3389.3900 ;
      RECT 3535.0800 3386.6900 3753.7200 3386.7900 ;
      RECT 3525.9200 3386.6900 3527.2200 3389.4900 ;
      RECT 3294.6200 3386.6900 3513.2600 3386.7900 ;
      RECT 3285.4600 3386.6900 3286.7600 3389.4900 ;
      RECT 3054.1600 3386.6900 3272.8000 3386.7900 ;
      RECT 3045.0000 3386.6900 3046.3000 3389.4900 ;
      RECT 2813.7000 3386.6900 3032.3400 3386.7900 ;
      RECT 2804.5400 3386.6900 2805.8400 3389.4900 ;
      RECT 2573.2400 3386.6900 2791.8800 3386.7900 ;
      RECT 2564.0800 3386.6900 2565.3800 3389.4900 ;
      RECT 2332.7800 3386.6900 2551.4200 3386.7900 ;
      RECT 2323.6200 3386.6900 2324.9200 3389.4900 ;
      RECT 2092.3200 3386.6900 2310.9600 3386.7900 ;
      RECT 2083.1600 3386.6900 2084.4600 3389.4900 ;
      RECT 1851.8600 3386.6900 2070.5000 3386.7900 ;
      RECT 1842.7000 3386.6900 1844.0000 3389.4900 ;
      RECT 1611.4000 3386.6900 1830.0400 3386.7900 ;
      RECT 1602.2400 3386.6900 1603.5400 3389.4900 ;
      RECT 1370.9400 3386.6900 1589.5800 3386.7900 ;
      RECT 1361.7800 3386.6900 1363.0800 3389.4900 ;
      RECT 1130.4800 3386.6900 1349.1200 3386.7900 ;
      RECT 1121.3200 3386.6900 1122.6200 3389.4900 ;
      RECT 890.0200 3386.6900 1108.6600 3386.7900 ;
      RECT 880.8600 3386.6900 882.1600 3389.4900 ;
      RECT 649.5600 3386.6900 868.2000 3386.7900 ;
      RECT 640.4000 3386.6900 641.7000 3389.4900 ;
      RECT 409.1000 3386.6900 627.7400 3386.7900 ;
      RECT 399.9400 3386.6900 401.2400 3389.4900 ;
      RECT 168.6400 3386.6900 387.2800 3386.7900 ;
      RECT 159.3800 3386.6900 160.6800 3389.4900 ;
      RECT 3776.3800 3382.8600 3777.7800 3387.6900 ;
      RECT 3770.3800 3382.8600 3773.7800 3617.3000 ;
      RECT 3816.2800 3380.8600 3817.6800 3390.1900 ;
      RECT 3780.3800 3380.8600 3813.6800 3387.6900 ;
      RECT 3756.3200 3380.8600 3763.7800 3393.8900 ;
      RECT 3529.9200 3380.8600 3753.7200 3386.6900 ;
      RECT 3515.8600 3380.8600 3523.3200 3393.8900 ;
      RECT 3289.4600 3380.8600 3513.2600 3386.6900 ;
      RECT 3275.4000 3380.8600 3282.8600 3393.8900 ;
      RECT 3049.0000 3380.8600 3272.8000 3386.6900 ;
      RECT 3034.9400 3380.8600 3042.4000 3393.8900 ;
      RECT 2808.5400 3380.8600 3032.3400 3386.6900 ;
      RECT 2794.4800 3380.8600 2801.9400 3393.8900 ;
      RECT 2568.0800 3380.8600 2791.8800 3386.6900 ;
      RECT 2554.0200 3380.8600 2561.4800 3393.8900 ;
      RECT 2327.6200 3380.8600 2551.4200 3386.6900 ;
      RECT 2313.5600 3380.8600 2321.0200 3393.8900 ;
      RECT 2087.1600 3380.8600 2310.9600 3386.6900 ;
      RECT 2073.1000 3380.8600 2080.5600 3393.8900 ;
      RECT 1846.7000 3380.8600 2070.5000 3386.6900 ;
      RECT 1832.6400 3380.8600 1840.1000 3393.8900 ;
      RECT 1606.2400 3380.8600 1830.0400 3386.6900 ;
      RECT 1592.1800 3380.8600 1599.6400 3393.8900 ;
      RECT 1365.7800 3380.8600 1589.5800 3386.6900 ;
      RECT 1351.7200 3380.8600 1359.1800 3393.8900 ;
      RECT 1125.3200 3380.8600 1349.1200 3386.6900 ;
      RECT 1111.2600 3380.8600 1118.7200 3393.8900 ;
      RECT 884.8600 3380.8600 1108.6600 3386.6900 ;
      RECT 870.8000 3380.8600 878.2600 3393.8900 ;
      RECT 644.4000 3380.8600 868.2000 3386.6900 ;
      RECT 630.3400 3380.8600 637.8000 3393.8900 ;
      RECT 403.9400 3380.8600 627.7400 3386.6900 ;
      RECT 389.8800 3380.8600 397.3400 3393.8900 ;
      RECT 163.3800 3380.8600 387.2800 3386.6900 ;
      RECT 3820.2800 3376.8600 3917.8400 3617.3000 ;
      RECT 3780.3800 3376.8600 3817.6800 3380.8600 ;
      RECT 3770.3800 3376.8600 3777.7800 3382.8600 ;
      RECT 3770.3800 3367.4600 3917.8400 3376.8600 ;
      RECT 3529.9200 3144.0500 3763.7800 3380.8600 ;
      RECT 3289.4600 3144.0500 3523.3200 3380.8600 ;
      RECT 3049.0000 3144.0500 3282.8600 3380.8600 ;
      RECT 2808.5400 3144.0500 3042.4000 3380.8600 ;
      RECT 2568.0800 3144.0500 2801.9400 3380.8600 ;
      RECT 2327.6200 3144.0500 2561.4800 3380.8600 ;
      RECT 2087.1600 3144.0500 2321.0200 3380.8600 ;
      RECT 1846.7000 3144.0500 2080.5600 3380.8600 ;
      RECT 1606.2400 3144.0500 1840.1000 3380.8600 ;
      RECT 1365.7800 3144.0500 1599.6400 3380.8600 ;
      RECT 1125.3200 3144.0500 1359.1800 3380.8600 ;
      RECT 884.8600 3144.0500 1118.7200 3380.8600 ;
      RECT 644.4000 3144.0500 878.2600 3380.8600 ;
      RECT 403.9400 3144.0500 637.8000 3380.8600 ;
      RECT 163.3800 3144.0500 397.3400 3380.8600 ;
      RECT 159.3800 3142.9100 160.7800 3386.6900 ;
      RECT 123.4800 3142.9100 156.7800 3388.0500 ;
      RECT 123.4800 3142.8100 150.4400 3142.9100 ;
      RECT 3816.2800 3142.6500 3817.6800 3367.4600 ;
      RECT 3780.3800 3142.6500 3813.6800 3367.4600 ;
      RECT 3780.3800 3142.5500 3807.3400 3142.6500 ;
      RECT 123.4800 3140.7100 149.7900 3142.8100 ;
      RECT 159.4800 3140.6100 160.7800 3142.9100 ;
      RECT 123.4800 3140.6100 150.4400 3140.7100 ;
      RECT 3780.3800 3140.4500 3806.6900 3142.5500 ;
      RECT 3816.3800 3140.3500 3817.6800 3142.6500 ;
      RECT 3780.3800 3140.3500 3807.3400 3140.4500 ;
      RECT 123.4800 3140.3100 156.7800 3140.6100 ;
      RECT 3780.3800 3140.1500 3813.6800 3140.3500 ;
      RECT 3776.3800 3140.1500 3777.7800 3367.4600 ;
      RECT 3784.2200 3140.0500 3813.6800 3140.1500 ;
      RECT 3529.9200 3139.6500 3753.7200 3144.0500 ;
      RECT 3525.9200 3139.6500 3527.3200 3386.6900 ;
      RECT 3289.4600 3139.6500 3513.2600 3144.0500 ;
      RECT 3285.4600 3139.6500 3286.8600 3386.6900 ;
      RECT 3049.0000 3139.6500 3272.8000 3144.0500 ;
      RECT 3045.0000 3139.6500 3046.4000 3386.6900 ;
      RECT 2808.5400 3139.6500 3032.3400 3144.0500 ;
      RECT 2804.5400 3139.6500 2805.9400 3386.6900 ;
      RECT 2568.0800 3139.6500 2791.8800 3144.0500 ;
      RECT 2564.0800 3139.6500 2565.4800 3386.6900 ;
      RECT 2327.6200 3139.6500 2551.4200 3144.0500 ;
      RECT 2323.6200 3139.6500 2325.0200 3386.6900 ;
      RECT 2087.1600 3139.6500 2310.9600 3144.0500 ;
      RECT 2083.1600 3139.6500 2084.5600 3386.6900 ;
      RECT 1846.7000 3139.6500 2070.5000 3144.0500 ;
      RECT 1842.7000 3139.6500 1844.1000 3386.6900 ;
      RECT 1606.2400 3139.6500 1830.0400 3144.0500 ;
      RECT 1602.2400 3139.6500 1603.6400 3386.6900 ;
      RECT 1365.7800 3139.6500 1589.5800 3144.0500 ;
      RECT 1361.7800 3139.6500 1363.1800 3386.6900 ;
      RECT 1125.3200 3139.6500 1349.1200 3144.0500 ;
      RECT 1121.3200 3139.6500 1122.7200 3386.6900 ;
      RECT 884.8600 3139.6500 1108.6600 3144.0500 ;
      RECT 880.8600 3139.6500 882.2600 3386.6900 ;
      RECT 644.4000 3139.6500 868.2000 3144.0500 ;
      RECT 640.4000 3139.6500 641.8000 3386.6900 ;
      RECT 403.9400 3139.6500 627.7400 3144.0500 ;
      RECT 399.9400 3139.6500 401.3400 3386.6900 ;
      RECT 163.3800 3139.6500 387.2800 3144.0500 ;
      RECT 159.3800 3139.6500 160.7800 3140.6100 ;
      RECT 3535.0800 3139.5500 3753.7200 3139.6500 ;
      RECT 3294.6200 3139.5500 3513.2600 3139.6500 ;
      RECT 3054.1600 3139.5500 3272.8000 3139.6500 ;
      RECT 2813.7000 3139.5500 3032.3400 3139.6500 ;
      RECT 2573.2400 3139.5500 2791.8800 3139.6500 ;
      RECT 2332.7800 3139.5500 2551.4200 3139.6500 ;
      RECT 2092.3200 3139.5500 2310.9600 3139.6500 ;
      RECT 1851.8600 3139.5500 2070.5000 3139.6500 ;
      RECT 1611.4000 3139.5500 1830.0400 3139.6500 ;
      RECT 1370.9400 3139.5500 1589.5800 3139.6500 ;
      RECT 1130.4800 3139.5500 1349.1200 3139.6500 ;
      RECT 890.0200 3139.5500 1108.6600 3139.6500 ;
      RECT 649.5600 3139.5500 868.2000 3139.6500 ;
      RECT 409.1000 3139.5500 627.7400 3139.6500 ;
      RECT 168.6400 3139.5500 387.2800 3139.6500 ;
      RECT 156.3100 3138.2100 156.7800 3140.3100 ;
      RECT 123.4800 3138.2100 151.7050 3140.3100 ;
      RECT 3784.8700 3137.9500 3813.6800 3140.0500 ;
      RECT 3784.2200 3137.8500 3813.6800 3137.9500 ;
      RECT 3776.3800 3137.8500 3777.6800 3140.1500 ;
      RECT 3536.4800 3136.9500 3753.7200 3139.5500 ;
      RECT 3296.0200 3136.9500 3513.2600 3139.5500 ;
      RECT 3055.5600 3136.9500 3272.8000 3139.5500 ;
      RECT 2815.1000 3136.9500 3032.3400 3139.5500 ;
      RECT 2574.6400 3136.9500 2791.8800 3139.5500 ;
      RECT 2334.1800 3136.9500 2551.4200 3139.5500 ;
      RECT 2093.7200 3136.9500 2310.9600 3139.5500 ;
      RECT 1853.2600 3136.9500 2070.5000 3139.5500 ;
      RECT 1612.8000 3136.9500 1830.0400 3139.5500 ;
      RECT 1372.3400 3136.9500 1589.5800 3139.5500 ;
      RECT 1131.8800 3136.9500 1349.1200 3139.5500 ;
      RECT 891.4200 3136.9500 1108.6600 3139.5500 ;
      RECT 650.9600 3136.9500 868.2000 3139.5500 ;
      RECT 410.5000 3136.9500 627.7400 3139.5500 ;
      RECT 170.0400 3136.9500 387.2800 3139.5500 ;
      RECT 3535.0800 3136.8500 3753.7200 3136.9500 ;
      RECT 3525.9200 3136.8500 3527.2200 3139.6500 ;
      RECT 3294.6200 3136.8500 3513.2600 3136.9500 ;
      RECT 3285.4600 3136.8500 3286.7600 3139.6500 ;
      RECT 3054.1600 3136.8500 3272.8000 3136.9500 ;
      RECT 3045.0000 3136.8500 3046.3000 3139.6500 ;
      RECT 2813.7000 3136.8500 3032.3400 3136.9500 ;
      RECT 2804.5400 3136.8500 2805.8400 3139.6500 ;
      RECT 2573.2400 3136.8500 2791.8800 3136.9500 ;
      RECT 2564.0800 3136.8500 2565.3800 3139.6500 ;
      RECT 2332.7800 3136.8500 2551.4200 3136.9500 ;
      RECT 2323.6200 3136.8500 2324.9200 3139.6500 ;
      RECT 2092.3200 3136.8500 2310.9600 3136.9500 ;
      RECT 2083.1600 3136.8500 2084.4600 3139.6500 ;
      RECT 1851.8600 3136.8500 2070.5000 3136.9500 ;
      RECT 1842.7000 3136.8500 1844.0000 3139.6500 ;
      RECT 1611.4000 3136.8500 1830.0400 3136.9500 ;
      RECT 1602.2400 3136.8500 1603.5400 3139.6500 ;
      RECT 1370.9400 3136.8500 1589.5800 3136.9500 ;
      RECT 1361.7800 3136.8500 1363.0800 3139.6500 ;
      RECT 1130.4800 3136.8500 1349.1200 3136.9500 ;
      RECT 1121.3200 3136.8500 1122.6200 3139.6500 ;
      RECT 890.0200 3136.8500 1108.6600 3136.9500 ;
      RECT 880.8600 3136.8500 882.1600 3139.6500 ;
      RECT 649.5600 3136.8500 868.2000 3136.9500 ;
      RECT 640.4000 3136.8500 641.7000 3139.6500 ;
      RECT 409.1000 3136.8500 627.7400 3136.9500 ;
      RECT 399.9400 3136.8500 401.2400 3139.6500 ;
      RECT 168.6400 3136.8500 387.2800 3136.9500 ;
      RECT 159.3800 3136.8500 160.6800 3139.6500 ;
      RECT 3776.3800 3133.0200 3777.7800 3137.8500 ;
      RECT 3770.3800 3133.0200 3773.7800 3367.4600 ;
      RECT 3816.2800 3131.0200 3817.6800 3140.3500 ;
      RECT 3780.3800 3131.0200 3813.6800 3137.8500 ;
      RECT 3756.3200 3131.0200 3763.7800 3144.0500 ;
      RECT 3529.9200 3131.0200 3753.7200 3136.8500 ;
      RECT 3515.8600 3131.0200 3523.3200 3144.0500 ;
      RECT 3289.4600 3131.0200 3513.2600 3136.8500 ;
      RECT 3275.4000 3131.0200 3282.8600 3144.0500 ;
      RECT 3049.0000 3131.0200 3272.8000 3136.8500 ;
      RECT 3034.9400 3131.0200 3042.4000 3144.0500 ;
      RECT 2808.5400 3131.0200 3032.3400 3136.8500 ;
      RECT 2794.4800 3131.0200 2801.9400 3144.0500 ;
      RECT 2568.0800 3131.0200 2791.8800 3136.8500 ;
      RECT 2554.0200 3131.0200 2561.4800 3144.0500 ;
      RECT 2327.6200 3131.0200 2551.4200 3136.8500 ;
      RECT 2313.5600 3131.0200 2321.0200 3144.0500 ;
      RECT 2087.1600 3131.0200 2310.9600 3136.8500 ;
      RECT 2073.1000 3131.0200 2080.5600 3144.0500 ;
      RECT 1846.7000 3131.0200 2070.5000 3136.8500 ;
      RECT 1832.6400 3131.0200 1840.1000 3144.0500 ;
      RECT 1606.2400 3131.0200 1830.0400 3136.8500 ;
      RECT 1592.1800 3131.0200 1599.6400 3144.0500 ;
      RECT 1365.7800 3131.0200 1589.5800 3136.8500 ;
      RECT 1351.7200 3131.0200 1359.1800 3144.0500 ;
      RECT 1125.3200 3131.0200 1349.1200 3136.8500 ;
      RECT 1111.2600 3131.0200 1118.7200 3144.0500 ;
      RECT 884.8600 3131.0200 1108.6600 3136.8500 ;
      RECT 870.8000 3131.0200 878.2600 3144.0500 ;
      RECT 644.4000 3131.0200 868.2000 3136.8500 ;
      RECT 630.3400 3131.0200 637.8000 3144.0500 ;
      RECT 403.9400 3131.0200 627.7400 3136.8500 ;
      RECT 389.8800 3131.0200 397.3400 3144.0500 ;
      RECT 163.3800 3131.0200 387.2800 3136.8500 ;
      RECT 3820.2800 3127.0200 3917.8400 3367.4600 ;
      RECT 3780.3800 3127.0200 3817.6800 3131.0200 ;
      RECT 3770.3800 3127.0200 3777.7800 3133.0200 ;
      RECT 3770.3800 3117.6200 3917.8400 3127.0200 ;
      RECT 3529.9200 2894.2100 3763.7800 3131.0200 ;
      RECT 3289.4600 2894.2100 3523.3200 3131.0200 ;
      RECT 3049.0000 2894.2100 3282.8600 3131.0200 ;
      RECT 2808.5400 2894.2100 3042.4000 3131.0200 ;
      RECT 2568.0800 2894.2100 2801.9400 3131.0200 ;
      RECT 2327.6200 2894.2100 2561.4800 3131.0200 ;
      RECT 2087.1600 2894.2100 2321.0200 3131.0200 ;
      RECT 1846.7000 2894.2100 2080.5600 3131.0200 ;
      RECT 1606.2400 2894.2100 1840.1000 3131.0200 ;
      RECT 1365.7800 2894.2100 1599.6400 3131.0200 ;
      RECT 1125.3200 2894.2100 1359.1800 3131.0200 ;
      RECT 884.8600 2894.2100 1118.7200 3131.0200 ;
      RECT 644.4000 2894.2100 878.2600 3131.0200 ;
      RECT 403.9400 2894.2100 637.8000 3131.0200 ;
      RECT 163.3800 2894.2100 397.3400 3131.0200 ;
      RECT 159.3800 2893.0700 160.7800 3136.8500 ;
      RECT 123.4800 2893.0700 156.7800 3138.2100 ;
      RECT 123.4800 2892.9700 150.4400 2893.0700 ;
      RECT 3816.2800 2892.8100 3817.6800 3117.6200 ;
      RECT 3780.3800 2892.8100 3813.6800 3117.6200 ;
      RECT 3780.3800 2892.7100 3807.3400 2892.8100 ;
      RECT 123.4800 2890.8700 149.7900 2892.9700 ;
      RECT 159.4800 2890.7700 160.7800 2893.0700 ;
      RECT 123.4800 2890.7700 150.4400 2890.8700 ;
      RECT 3780.3800 2890.6100 3806.6900 2892.7100 ;
      RECT 3816.3800 2890.5100 3817.6800 2892.8100 ;
      RECT 3780.3800 2890.5100 3807.3400 2890.6100 ;
      RECT 123.4800 2890.4700 156.7800 2890.7700 ;
      RECT 3780.3800 2890.3100 3813.6800 2890.5100 ;
      RECT 3776.3800 2890.3100 3777.7800 3117.6200 ;
      RECT 3784.2200 2890.2100 3813.6800 2890.3100 ;
      RECT 3529.9200 2889.8100 3753.7200 2894.2100 ;
      RECT 3525.9200 2889.8100 3527.3200 3136.8500 ;
      RECT 3289.4600 2889.8100 3513.2600 2894.2100 ;
      RECT 3285.4600 2889.8100 3286.8600 3136.8500 ;
      RECT 3049.0000 2889.8100 3272.8000 2894.2100 ;
      RECT 3045.0000 2889.8100 3046.4000 3136.8500 ;
      RECT 2808.5400 2889.8100 3032.3400 2894.2100 ;
      RECT 2804.5400 2889.8100 2805.9400 3136.8500 ;
      RECT 2568.0800 2889.8100 2791.8800 2894.2100 ;
      RECT 2564.0800 2889.8100 2565.4800 3136.8500 ;
      RECT 2327.6200 2889.8100 2551.4200 2894.2100 ;
      RECT 2323.6200 2889.8100 2325.0200 3136.8500 ;
      RECT 2087.1600 2889.8100 2310.9600 2894.2100 ;
      RECT 2083.1600 2889.8100 2084.5600 3136.8500 ;
      RECT 1846.7000 2889.8100 2070.5000 2894.2100 ;
      RECT 1842.7000 2889.8100 1844.1000 3136.8500 ;
      RECT 1606.2400 2889.8100 1830.0400 2894.2100 ;
      RECT 1602.2400 2889.8100 1603.6400 3136.8500 ;
      RECT 1365.7800 2889.8100 1589.5800 2894.2100 ;
      RECT 1361.7800 2889.8100 1363.1800 3136.8500 ;
      RECT 1125.3200 2889.8100 1349.1200 2894.2100 ;
      RECT 1121.3200 2889.8100 1122.7200 3136.8500 ;
      RECT 884.8600 2889.8100 1108.6600 2894.2100 ;
      RECT 880.8600 2889.8100 882.2600 3136.8500 ;
      RECT 644.4000 2889.8100 868.2000 2894.2100 ;
      RECT 640.4000 2889.8100 641.8000 3136.8500 ;
      RECT 403.9400 2889.8100 627.7400 2894.2100 ;
      RECT 399.9400 2889.8100 401.3400 3136.8500 ;
      RECT 163.3800 2889.8100 387.2800 2894.2100 ;
      RECT 159.3800 2889.8100 160.7800 2890.7700 ;
      RECT 3535.0800 2889.7100 3753.7200 2889.8100 ;
      RECT 3294.6200 2889.7100 3513.2600 2889.8100 ;
      RECT 3054.1600 2889.7100 3272.8000 2889.8100 ;
      RECT 2813.7000 2889.7100 3032.3400 2889.8100 ;
      RECT 2573.2400 2889.7100 2791.8800 2889.8100 ;
      RECT 2332.7800 2889.7100 2551.4200 2889.8100 ;
      RECT 2092.3200 2889.7100 2310.9600 2889.8100 ;
      RECT 1851.8600 2889.7100 2070.5000 2889.8100 ;
      RECT 1611.4000 2889.7100 1830.0400 2889.8100 ;
      RECT 1370.9400 2889.7100 1589.5800 2889.8100 ;
      RECT 1130.4800 2889.7100 1349.1200 2889.8100 ;
      RECT 890.0200 2889.7100 1108.6600 2889.8100 ;
      RECT 649.5600 2889.7100 868.2000 2889.8100 ;
      RECT 409.1000 2889.7100 627.7400 2889.8100 ;
      RECT 168.6400 2889.7100 387.2800 2889.8100 ;
      RECT 156.3100 2888.3700 156.7800 2890.4700 ;
      RECT 123.4800 2888.3700 151.7050 2890.4700 ;
      RECT 3784.8700 2888.1100 3813.6800 2890.2100 ;
      RECT 3784.2200 2888.0100 3813.6800 2888.1100 ;
      RECT 3776.3800 2888.0100 3777.6800 2890.3100 ;
      RECT 3536.4800 2887.1100 3753.7200 2889.7100 ;
      RECT 3296.0200 2887.1100 3513.2600 2889.7100 ;
      RECT 3055.5600 2887.1100 3272.8000 2889.7100 ;
      RECT 2815.1000 2887.1100 3032.3400 2889.7100 ;
      RECT 2574.6400 2887.1100 2791.8800 2889.7100 ;
      RECT 2334.1800 2887.1100 2551.4200 2889.7100 ;
      RECT 2093.7200 2887.1100 2310.9600 2889.7100 ;
      RECT 1853.2600 2887.1100 2070.5000 2889.7100 ;
      RECT 1612.8000 2887.1100 1830.0400 2889.7100 ;
      RECT 1372.3400 2887.1100 1589.5800 2889.7100 ;
      RECT 1131.8800 2887.1100 1349.1200 2889.7100 ;
      RECT 891.4200 2887.1100 1108.6600 2889.7100 ;
      RECT 650.9600 2887.1100 868.2000 2889.7100 ;
      RECT 410.5000 2887.1100 627.7400 2889.7100 ;
      RECT 170.0400 2887.1100 387.2800 2889.7100 ;
      RECT 3535.0800 2887.0100 3753.7200 2887.1100 ;
      RECT 3525.9200 2887.0100 3527.2200 2889.8100 ;
      RECT 3294.6200 2887.0100 3513.2600 2887.1100 ;
      RECT 3285.4600 2887.0100 3286.7600 2889.8100 ;
      RECT 3054.1600 2887.0100 3272.8000 2887.1100 ;
      RECT 3045.0000 2887.0100 3046.3000 2889.8100 ;
      RECT 2813.7000 2887.0100 3032.3400 2887.1100 ;
      RECT 2804.5400 2887.0100 2805.8400 2889.8100 ;
      RECT 2573.2400 2887.0100 2791.8800 2887.1100 ;
      RECT 2564.0800 2887.0100 2565.3800 2889.8100 ;
      RECT 2332.7800 2887.0100 2551.4200 2887.1100 ;
      RECT 2323.6200 2887.0100 2324.9200 2889.8100 ;
      RECT 2092.3200 2887.0100 2310.9600 2887.1100 ;
      RECT 2083.1600 2887.0100 2084.4600 2889.8100 ;
      RECT 1851.8600 2887.0100 2070.5000 2887.1100 ;
      RECT 1842.7000 2887.0100 1844.0000 2889.8100 ;
      RECT 1611.4000 2887.0100 1830.0400 2887.1100 ;
      RECT 1602.2400 2887.0100 1603.5400 2889.8100 ;
      RECT 1370.9400 2887.0100 1589.5800 2887.1100 ;
      RECT 1361.7800 2887.0100 1363.0800 2889.8100 ;
      RECT 1130.4800 2887.0100 1349.1200 2887.1100 ;
      RECT 1121.3200 2887.0100 1122.6200 2889.8100 ;
      RECT 890.0200 2887.0100 1108.6600 2887.1100 ;
      RECT 880.8600 2887.0100 882.1600 2889.8100 ;
      RECT 649.5600 2887.0100 868.2000 2887.1100 ;
      RECT 640.4000 2887.0100 641.7000 2889.8100 ;
      RECT 409.1000 2887.0100 627.7400 2887.1100 ;
      RECT 399.9400 2887.0100 401.2400 2889.8100 ;
      RECT 168.6400 2887.0100 387.2800 2887.1100 ;
      RECT 159.3800 2887.0100 160.6800 2889.8100 ;
      RECT 3776.3800 2883.1800 3777.7800 2888.0100 ;
      RECT 3770.3800 2883.1800 3773.7800 3117.6200 ;
      RECT 3816.2800 2881.1800 3817.6800 2890.5100 ;
      RECT 3780.3800 2881.1800 3813.6800 2888.0100 ;
      RECT 3756.3200 2881.1800 3763.7800 2894.2100 ;
      RECT 3529.9200 2881.1800 3753.7200 2887.0100 ;
      RECT 3515.8600 2881.1800 3523.3200 2894.2100 ;
      RECT 3289.4600 2881.1800 3513.2600 2887.0100 ;
      RECT 3275.4000 2881.1800 3282.8600 2894.2100 ;
      RECT 3049.0000 2881.1800 3272.8000 2887.0100 ;
      RECT 3034.9400 2881.1800 3042.4000 2894.2100 ;
      RECT 2808.5400 2881.1800 3032.3400 2887.0100 ;
      RECT 2794.4800 2881.1800 2801.9400 2894.2100 ;
      RECT 2568.0800 2881.1800 2791.8800 2887.0100 ;
      RECT 2554.0200 2881.1800 2561.4800 2894.2100 ;
      RECT 2327.6200 2881.1800 2551.4200 2887.0100 ;
      RECT 2313.5600 2881.1800 2321.0200 2894.2100 ;
      RECT 2087.1600 2881.1800 2310.9600 2887.0100 ;
      RECT 2073.1000 2881.1800 2080.5600 2894.2100 ;
      RECT 1846.7000 2881.1800 2070.5000 2887.0100 ;
      RECT 1832.6400 2881.1800 1840.1000 2894.2100 ;
      RECT 1606.2400 2881.1800 1830.0400 2887.0100 ;
      RECT 1592.1800 2881.1800 1599.6400 2894.2100 ;
      RECT 1365.7800 2881.1800 1589.5800 2887.0100 ;
      RECT 1351.7200 2881.1800 1359.1800 2894.2100 ;
      RECT 1125.3200 2881.1800 1349.1200 2887.0100 ;
      RECT 1111.2600 2881.1800 1118.7200 2894.2100 ;
      RECT 884.8600 2881.1800 1108.6600 2887.0100 ;
      RECT 870.8000 2881.1800 878.2600 2894.2100 ;
      RECT 644.4000 2881.1800 868.2000 2887.0100 ;
      RECT 630.3400 2881.1800 637.8000 2894.2100 ;
      RECT 403.9400 2881.1800 627.7400 2887.0100 ;
      RECT 389.8800 2881.1800 397.3400 2894.2100 ;
      RECT 163.3800 2881.1800 387.2800 2887.0100 ;
      RECT 3820.2800 2877.1800 3917.8400 3117.6200 ;
      RECT 3780.3800 2877.1800 3817.6800 2881.1800 ;
      RECT 3770.3800 2877.1800 3777.7800 2883.1800 ;
      RECT 3770.3800 2867.7800 3917.8400 2877.1800 ;
      RECT 3529.9200 2644.3700 3763.7800 2881.1800 ;
      RECT 3289.4600 2644.3700 3523.3200 2881.1800 ;
      RECT 3049.0000 2644.3700 3282.8600 2881.1800 ;
      RECT 2808.5400 2644.3700 3042.4000 2881.1800 ;
      RECT 2568.0800 2644.3700 2801.9400 2881.1800 ;
      RECT 2327.6200 2644.3700 2561.4800 2881.1800 ;
      RECT 2087.1600 2644.3700 2321.0200 2881.1800 ;
      RECT 1846.7000 2644.3700 2080.5600 2881.1800 ;
      RECT 1606.2400 2644.3700 1840.1000 2881.1800 ;
      RECT 1365.7800 2644.3700 1599.6400 2881.1800 ;
      RECT 1125.3200 2644.3700 1359.1800 2881.1800 ;
      RECT 884.8600 2644.3700 1118.7200 2881.1800 ;
      RECT 644.4000 2644.3700 878.2600 2881.1800 ;
      RECT 403.9400 2644.3700 637.8000 2881.1800 ;
      RECT 163.3800 2644.3700 397.3400 2881.1800 ;
      RECT 159.3800 2643.2300 160.7800 2887.0100 ;
      RECT 123.4800 2643.2300 156.7800 2888.3700 ;
      RECT 123.4800 2643.1300 150.4400 2643.2300 ;
      RECT 3816.2800 2642.9700 3817.6800 2867.7800 ;
      RECT 3780.3800 2642.9700 3813.6800 2867.7800 ;
      RECT 3780.3800 2642.8700 3807.3400 2642.9700 ;
      RECT 123.4800 2641.0300 149.7900 2643.1300 ;
      RECT 159.4800 2640.9300 160.7800 2643.2300 ;
      RECT 123.4800 2640.9300 150.4400 2641.0300 ;
      RECT 3780.3800 2640.7700 3806.6900 2642.8700 ;
      RECT 3816.3800 2640.6700 3817.6800 2642.9700 ;
      RECT 3780.3800 2640.6700 3807.3400 2640.7700 ;
      RECT 123.4800 2640.6300 156.7800 2640.9300 ;
      RECT 3780.3800 2640.4700 3813.6800 2640.6700 ;
      RECT 3776.3800 2640.4700 3777.7800 2867.7800 ;
      RECT 3784.2200 2640.3700 3813.6800 2640.4700 ;
      RECT 3529.9200 2639.9700 3753.7200 2644.3700 ;
      RECT 3525.9200 2639.9700 3527.3200 2887.0100 ;
      RECT 3289.4600 2639.9700 3513.2600 2644.3700 ;
      RECT 3285.4600 2639.9700 3286.8600 2887.0100 ;
      RECT 3049.0000 2639.9700 3272.8000 2644.3700 ;
      RECT 3045.0000 2639.9700 3046.4000 2887.0100 ;
      RECT 2808.5400 2639.9700 3032.3400 2644.3700 ;
      RECT 2804.5400 2639.9700 2805.9400 2887.0100 ;
      RECT 2568.0800 2639.9700 2791.8800 2644.3700 ;
      RECT 2564.0800 2639.9700 2565.4800 2887.0100 ;
      RECT 2327.6200 2639.9700 2551.4200 2644.3700 ;
      RECT 2323.6200 2639.9700 2325.0200 2887.0100 ;
      RECT 2087.1600 2639.9700 2310.9600 2644.3700 ;
      RECT 2083.1600 2639.9700 2084.5600 2887.0100 ;
      RECT 1846.7000 2639.9700 2070.5000 2644.3700 ;
      RECT 1842.7000 2639.9700 1844.1000 2887.0100 ;
      RECT 1606.2400 2639.9700 1830.0400 2644.3700 ;
      RECT 1602.2400 2639.9700 1603.6400 2887.0100 ;
      RECT 1365.7800 2639.9700 1589.5800 2644.3700 ;
      RECT 1361.7800 2639.9700 1363.1800 2887.0100 ;
      RECT 1125.3200 2639.9700 1349.1200 2644.3700 ;
      RECT 1121.3200 2639.9700 1122.7200 2887.0100 ;
      RECT 884.8600 2639.9700 1108.6600 2644.3700 ;
      RECT 880.8600 2639.9700 882.2600 2887.0100 ;
      RECT 644.4000 2639.9700 868.2000 2644.3700 ;
      RECT 640.4000 2639.9700 641.8000 2887.0100 ;
      RECT 403.9400 2639.9700 627.7400 2644.3700 ;
      RECT 399.9400 2639.9700 401.3400 2887.0100 ;
      RECT 163.3800 2639.9700 387.2800 2644.3700 ;
      RECT 159.3800 2639.9700 160.7800 2640.9300 ;
      RECT 3535.0800 2639.8700 3753.7200 2639.9700 ;
      RECT 3294.6200 2639.8700 3513.2600 2639.9700 ;
      RECT 3054.1600 2639.8700 3272.8000 2639.9700 ;
      RECT 2813.7000 2639.8700 3032.3400 2639.9700 ;
      RECT 2573.2400 2639.8700 2791.8800 2639.9700 ;
      RECT 2332.7800 2639.8700 2551.4200 2639.9700 ;
      RECT 2092.3200 2639.8700 2310.9600 2639.9700 ;
      RECT 1851.8600 2639.8700 2070.5000 2639.9700 ;
      RECT 1611.4000 2639.8700 1830.0400 2639.9700 ;
      RECT 1370.9400 2639.8700 1589.5800 2639.9700 ;
      RECT 1130.4800 2639.8700 1349.1200 2639.9700 ;
      RECT 890.0200 2639.8700 1108.6600 2639.9700 ;
      RECT 649.5600 2639.8700 868.2000 2639.9700 ;
      RECT 409.1000 2639.8700 627.7400 2639.9700 ;
      RECT 168.6400 2639.8700 387.2800 2639.9700 ;
      RECT 156.3100 2638.5300 156.7800 2640.6300 ;
      RECT 123.4800 2638.5300 151.7050 2640.6300 ;
      RECT 3784.8700 2638.2700 3813.6800 2640.3700 ;
      RECT 3784.2200 2638.1700 3813.6800 2638.2700 ;
      RECT 3776.3800 2638.1700 3777.6800 2640.4700 ;
      RECT 3536.4800 2637.2700 3753.7200 2639.8700 ;
      RECT 3296.0200 2637.2700 3513.2600 2639.8700 ;
      RECT 3055.5600 2637.2700 3272.8000 2639.8700 ;
      RECT 2815.1000 2637.2700 3032.3400 2639.8700 ;
      RECT 2574.6400 2637.2700 2791.8800 2639.8700 ;
      RECT 2334.1800 2637.2700 2551.4200 2639.8700 ;
      RECT 2093.7200 2637.2700 2310.9600 2639.8700 ;
      RECT 1853.2600 2637.2700 2070.5000 2639.8700 ;
      RECT 1612.8000 2637.2700 1830.0400 2639.8700 ;
      RECT 1372.3400 2637.2700 1589.5800 2639.8700 ;
      RECT 1131.8800 2637.2700 1349.1200 2639.8700 ;
      RECT 891.4200 2637.2700 1108.6600 2639.8700 ;
      RECT 650.9600 2637.2700 868.2000 2639.8700 ;
      RECT 410.5000 2637.2700 627.7400 2639.8700 ;
      RECT 170.0400 2637.2700 387.2800 2639.8700 ;
      RECT 3535.0800 2637.1700 3753.7200 2637.2700 ;
      RECT 3525.9200 2637.1700 3527.2200 2639.9700 ;
      RECT 3294.6200 2637.1700 3513.2600 2637.2700 ;
      RECT 3285.4600 2637.1700 3286.7600 2639.9700 ;
      RECT 3054.1600 2637.1700 3272.8000 2637.2700 ;
      RECT 3045.0000 2637.1700 3046.3000 2639.9700 ;
      RECT 2813.7000 2637.1700 3032.3400 2637.2700 ;
      RECT 2804.5400 2637.1700 2805.8400 2639.9700 ;
      RECT 2573.2400 2637.1700 2791.8800 2637.2700 ;
      RECT 2564.0800 2637.1700 2565.3800 2639.9700 ;
      RECT 2332.7800 2637.1700 2551.4200 2637.2700 ;
      RECT 2323.6200 2637.1700 2324.9200 2639.9700 ;
      RECT 2092.3200 2637.1700 2310.9600 2637.2700 ;
      RECT 2083.1600 2637.1700 2084.4600 2639.9700 ;
      RECT 1851.8600 2637.1700 2070.5000 2637.2700 ;
      RECT 1842.7000 2637.1700 1844.0000 2639.9700 ;
      RECT 1611.4000 2637.1700 1830.0400 2637.2700 ;
      RECT 1602.2400 2637.1700 1603.5400 2639.9700 ;
      RECT 1370.9400 2637.1700 1589.5800 2637.2700 ;
      RECT 1361.7800 2637.1700 1363.0800 2639.9700 ;
      RECT 1130.4800 2637.1700 1349.1200 2637.2700 ;
      RECT 1121.3200 2637.1700 1122.6200 2639.9700 ;
      RECT 890.0200 2637.1700 1108.6600 2637.2700 ;
      RECT 880.8600 2637.1700 882.1600 2639.9700 ;
      RECT 649.5600 2637.1700 868.2000 2637.2700 ;
      RECT 640.4000 2637.1700 641.7000 2639.9700 ;
      RECT 409.1000 2637.1700 627.7400 2637.2700 ;
      RECT 399.9400 2637.1700 401.2400 2639.9700 ;
      RECT 168.6400 2637.1700 387.2800 2637.2700 ;
      RECT 159.3800 2637.1700 160.6800 2639.9700 ;
      RECT 3776.3800 2633.3400 3777.7800 2638.1700 ;
      RECT 3770.3800 2633.3400 3773.7800 2867.7800 ;
      RECT 3816.2800 2631.3400 3817.6800 2640.6700 ;
      RECT 3780.3800 2631.3400 3813.6800 2638.1700 ;
      RECT 3756.3200 2631.3400 3763.7800 2644.3700 ;
      RECT 3529.9200 2631.3400 3753.7200 2637.1700 ;
      RECT 3515.8600 2631.3400 3523.3200 2644.3700 ;
      RECT 3289.4600 2631.3400 3513.2600 2637.1700 ;
      RECT 3275.4000 2631.3400 3282.8600 2644.3700 ;
      RECT 3049.0000 2631.3400 3272.8000 2637.1700 ;
      RECT 3034.9400 2631.3400 3042.4000 2644.3700 ;
      RECT 2808.5400 2631.3400 3032.3400 2637.1700 ;
      RECT 2794.4800 2631.3400 2801.9400 2644.3700 ;
      RECT 2568.0800 2631.3400 2791.8800 2637.1700 ;
      RECT 2554.0200 2631.3400 2561.4800 2644.3700 ;
      RECT 2327.6200 2631.3400 2551.4200 2637.1700 ;
      RECT 2313.5600 2631.3400 2321.0200 2644.3700 ;
      RECT 2087.1600 2631.3400 2310.9600 2637.1700 ;
      RECT 2073.1000 2631.3400 2080.5600 2644.3700 ;
      RECT 1846.7000 2631.3400 2070.5000 2637.1700 ;
      RECT 1832.6400 2631.3400 1840.1000 2644.3700 ;
      RECT 1606.2400 2631.3400 1830.0400 2637.1700 ;
      RECT 1592.1800 2631.3400 1599.6400 2644.3700 ;
      RECT 1365.7800 2631.3400 1589.5800 2637.1700 ;
      RECT 1351.7200 2631.3400 1359.1800 2644.3700 ;
      RECT 1125.3200 2631.3400 1349.1200 2637.1700 ;
      RECT 1111.2600 2631.3400 1118.7200 2644.3700 ;
      RECT 884.8600 2631.3400 1108.6600 2637.1700 ;
      RECT 870.8000 2631.3400 878.2600 2644.3700 ;
      RECT 644.4000 2631.3400 868.2000 2637.1700 ;
      RECT 630.3400 2631.3400 637.8000 2644.3700 ;
      RECT 403.9400 2631.3400 627.7400 2637.1700 ;
      RECT 389.8800 2631.3400 397.3400 2644.3700 ;
      RECT 163.3800 2631.3400 387.2800 2637.1700 ;
      RECT 3820.2800 2627.3400 3917.8400 2867.7800 ;
      RECT 3780.3800 2627.3400 3817.6800 2631.3400 ;
      RECT 3770.3800 2627.3400 3777.7800 2633.3400 ;
      RECT 3770.3800 2617.9400 3917.8400 2627.3400 ;
      RECT 3529.9200 2394.5300 3763.7800 2631.3400 ;
      RECT 3289.4600 2394.5300 3523.3200 2631.3400 ;
      RECT 3049.0000 2394.5300 3282.8600 2631.3400 ;
      RECT 2808.5400 2394.5300 3042.4000 2631.3400 ;
      RECT 2568.0800 2394.5300 2801.9400 2631.3400 ;
      RECT 2327.6200 2394.5300 2561.4800 2631.3400 ;
      RECT 2087.1600 2394.5300 2321.0200 2631.3400 ;
      RECT 1846.7000 2394.5300 2080.5600 2631.3400 ;
      RECT 1606.2400 2394.5300 1840.1000 2631.3400 ;
      RECT 1365.7800 2394.5300 1599.6400 2631.3400 ;
      RECT 1125.3200 2394.5300 1359.1800 2631.3400 ;
      RECT 884.8600 2394.5300 1118.7200 2631.3400 ;
      RECT 644.4000 2394.5300 878.2600 2631.3400 ;
      RECT 403.9400 2394.5300 637.8000 2631.3400 ;
      RECT 163.3800 2394.5300 397.3400 2631.3400 ;
      RECT 159.3800 2393.3900 160.7800 2637.1700 ;
      RECT 123.4800 2393.3900 156.7800 2638.5300 ;
      RECT 123.4800 2393.2900 150.4400 2393.3900 ;
      RECT 3816.2800 2393.1300 3817.6800 2617.9400 ;
      RECT 3780.3800 2393.1300 3813.6800 2617.9400 ;
      RECT 3780.3800 2393.0300 3807.3400 2393.1300 ;
      RECT 123.4800 2391.1900 149.7900 2393.2900 ;
      RECT 159.4800 2391.0900 160.7800 2393.3900 ;
      RECT 123.4800 2391.0900 150.4400 2391.1900 ;
      RECT 3780.3800 2390.9300 3806.6900 2393.0300 ;
      RECT 3816.3800 2390.8300 3817.6800 2393.1300 ;
      RECT 3780.3800 2390.8300 3807.3400 2390.9300 ;
      RECT 123.4800 2390.7900 156.7800 2391.0900 ;
      RECT 3780.3800 2390.6300 3813.6800 2390.8300 ;
      RECT 3776.3800 2390.6300 3777.7800 2617.9400 ;
      RECT 3784.2200 2390.5300 3813.6800 2390.6300 ;
      RECT 3529.9200 2390.1300 3753.7200 2394.5300 ;
      RECT 3525.9200 2390.1300 3527.3200 2637.1700 ;
      RECT 3289.4600 2390.1300 3513.2600 2394.5300 ;
      RECT 3285.4600 2390.1300 3286.8600 2637.1700 ;
      RECT 3049.0000 2390.1300 3272.8000 2394.5300 ;
      RECT 3045.0000 2390.1300 3046.4000 2637.1700 ;
      RECT 2808.5400 2390.1300 3032.3400 2394.5300 ;
      RECT 2804.5400 2390.1300 2805.9400 2637.1700 ;
      RECT 2568.0800 2390.1300 2791.8800 2394.5300 ;
      RECT 2564.0800 2390.1300 2565.4800 2637.1700 ;
      RECT 2327.6200 2390.1300 2551.4200 2394.5300 ;
      RECT 2323.6200 2390.1300 2325.0200 2637.1700 ;
      RECT 2087.1600 2390.1300 2310.9600 2394.5300 ;
      RECT 2083.1600 2390.1300 2084.5600 2637.1700 ;
      RECT 1846.7000 2390.1300 2070.5000 2394.5300 ;
      RECT 1842.7000 2390.1300 1844.1000 2637.1700 ;
      RECT 1606.2400 2390.1300 1830.0400 2394.5300 ;
      RECT 1602.2400 2390.1300 1603.6400 2637.1700 ;
      RECT 1365.7800 2390.1300 1589.5800 2394.5300 ;
      RECT 1361.7800 2390.1300 1363.1800 2637.1700 ;
      RECT 1125.3200 2390.1300 1349.1200 2394.5300 ;
      RECT 1121.3200 2390.1300 1122.7200 2637.1700 ;
      RECT 884.8600 2390.1300 1108.6600 2394.5300 ;
      RECT 880.8600 2390.1300 882.2600 2637.1700 ;
      RECT 644.4000 2390.1300 868.2000 2394.5300 ;
      RECT 640.4000 2390.1300 641.8000 2637.1700 ;
      RECT 403.9400 2390.1300 627.7400 2394.5300 ;
      RECT 399.9400 2390.1300 401.3400 2637.1700 ;
      RECT 163.3800 2390.1300 387.2800 2394.5300 ;
      RECT 159.3800 2390.1300 160.7800 2391.0900 ;
      RECT 3535.0800 2390.0300 3753.7200 2390.1300 ;
      RECT 3294.6200 2390.0300 3513.2600 2390.1300 ;
      RECT 3054.1600 2390.0300 3272.8000 2390.1300 ;
      RECT 2813.7000 2390.0300 3032.3400 2390.1300 ;
      RECT 2573.2400 2390.0300 2791.8800 2390.1300 ;
      RECT 2332.7800 2390.0300 2551.4200 2390.1300 ;
      RECT 2092.3200 2390.0300 2310.9600 2390.1300 ;
      RECT 1851.8600 2390.0300 2070.5000 2390.1300 ;
      RECT 1611.4000 2390.0300 1830.0400 2390.1300 ;
      RECT 1370.9400 2390.0300 1589.5800 2390.1300 ;
      RECT 1130.4800 2390.0300 1349.1200 2390.1300 ;
      RECT 890.0200 2390.0300 1108.6600 2390.1300 ;
      RECT 649.5600 2390.0300 868.2000 2390.1300 ;
      RECT 409.1000 2390.0300 627.7400 2390.1300 ;
      RECT 168.6400 2390.0300 387.2800 2390.1300 ;
      RECT 156.3100 2388.6900 156.7800 2390.7900 ;
      RECT 123.4800 2388.6900 151.7050 2390.7900 ;
      RECT 3784.8700 2388.4300 3813.6800 2390.5300 ;
      RECT 3784.2200 2388.3300 3813.6800 2388.4300 ;
      RECT 3776.3800 2388.3300 3777.6800 2390.6300 ;
      RECT 3536.4800 2387.4300 3753.7200 2390.0300 ;
      RECT 3296.0200 2387.4300 3513.2600 2390.0300 ;
      RECT 3055.5600 2387.4300 3272.8000 2390.0300 ;
      RECT 2815.1000 2387.4300 3032.3400 2390.0300 ;
      RECT 2574.6400 2387.4300 2791.8800 2390.0300 ;
      RECT 2334.1800 2387.4300 2551.4200 2390.0300 ;
      RECT 2093.7200 2387.4300 2310.9600 2390.0300 ;
      RECT 1853.2600 2387.4300 2070.5000 2390.0300 ;
      RECT 1612.8000 2387.4300 1830.0400 2390.0300 ;
      RECT 1372.3400 2387.4300 1589.5800 2390.0300 ;
      RECT 1131.8800 2387.4300 1349.1200 2390.0300 ;
      RECT 891.4200 2387.4300 1108.6600 2390.0300 ;
      RECT 650.9600 2387.4300 868.2000 2390.0300 ;
      RECT 410.5000 2387.4300 627.7400 2390.0300 ;
      RECT 170.0400 2387.4300 387.2800 2390.0300 ;
      RECT 3535.0800 2387.3300 3753.7200 2387.4300 ;
      RECT 3525.9200 2387.3300 3527.2200 2390.1300 ;
      RECT 3294.6200 2387.3300 3513.2600 2387.4300 ;
      RECT 3285.4600 2387.3300 3286.7600 2390.1300 ;
      RECT 3054.1600 2387.3300 3272.8000 2387.4300 ;
      RECT 3045.0000 2387.3300 3046.3000 2390.1300 ;
      RECT 2813.7000 2387.3300 3032.3400 2387.4300 ;
      RECT 2804.5400 2387.3300 2805.8400 2390.1300 ;
      RECT 2573.2400 2387.3300 2791.8800 2387.4300 ;
      RECT 2564.0800 2387.3300 2565.3800 2390.1300 ;
      RECT 2332.7800 2387.3300 2551.4200 2387.4300 ;
      RECT 2323.6200 2387.3300 2324.9200 2390.1300 ;
      RECT 2092.3200 2387.3300 2310.9600 2387.4300 ;
      RECT 2083.1600 2387.3300 2084.4600 2390.1300 ;
      RECT 1851.8600 2387.3300 2070.5000 2387.4300 ;
      RECT 1842.7000 2387.3300 1844.0000 2390.1300 ;
      RECT 1611.4000 2387.3300 1830.0400 2387.4300 ;
      RECT 1602.2400 2387.3300 1603.5400 2390.1300 ;
      RECT 1370.9400 2387.3300 1589.5800 2387.4300 ;
      RECT 1361.7800 2387.3300 1363.0800 2390.1300 ;
      RECT 1130.4800 2387.3300 1349.1200 2387.4300 ;
      RECT 1121.3200 2387.3300 1122.6200 2390.1300 ;
      RECT 890.0200 2387.3300 1108.6600 2387.4300 ;
      RECT 880.8600 2387.3300 882.1600 2390.1300 ;
      RECT 649.5600 2387.3300 868.2000 2387.4300 ;
      RECT 640.4000 2387.3300 641.7000 2390.1300 ;
      RECT 409.1000 2387.3300 627.7400 2387.4300 ;
      RECT 399.9400 2387.3300 401.2400 2390.1300 ;
      RECT 168.6400 2387.3300 387.2800 2387.4300 ;
      RECT 159.3800 2387.3300 160.6800 2390.1300 ;
      RECT 3776.3800 2383.5000 3777.7800 2388.3300 ;
      RECT 3770.3800 2383.5000 3773.7800 2617.9400 ;
      RECT 3816.2800 2381.5000 3817.6800 2390.8300 ;
      RECT 3780.3800 2381.5000 3813.6800 2388.3300 ;
      RECT 3756.3200 2381.5000 3763.7800 2394.5300 ;
      RECT 3529.9200 2381.5000 3753.7200 2387.3300 ;
      RECT 3515.8600 2381.5000 3523.3200 2394.5300 ;
      RECT 3289.4600 2381.5000 3513.2600 2387.3300 ;
      RECT 3275.4000 2381.5000 3282.8600 2394.5300 ;
      RECT 3049.0000 2381.5000 3272.8000 2387.3300 ;
      RECT 3034.9400 2381.5000 3042.4000 2394.5300 ;
      RECT 2808.5400 2381.5000 3032.3400 2387.3300 ;
      RECT 2794.4800 2381.5000 2801.9400 2394.5300 ;
      RECT 2568.0800 2381.5000 2791.8800 2387.3300 ;
      RECT 2554.0200 2381.5000 2561.4800 2394.5300 ;
      RECT 2327.6200 2381.5000 2551.4200 2387.3300 ;
      RECT 2313.5600 2381.5000 2321.0200 2394.5300 ;
      RECT 2087.1600 2381.5000 2310.9600 2387.3300 ;
      RECT 2073.1000 2381.5000 2080.5600 2394.5300 ;
      RECT 1846.7000 2381.5000 2070.5000 2387.3300 ;
      RECT 1832.6400 2381.5000 1840.1000 2394.5300 ;
      RECT 1606.2400 2381.5000 1830.0400 2387.3300 ;
      RECT 1592.1800 2381.5000 1599.6400 2394.5300 ;
      RECT 1365.7800 2381.5000 1589.5800 2387.3300 ;
      RECT 1351.7200 2381.5000 1359.1800 2394.5300 ;
      RECT 1125.3200 2381.5000 1349.1200 2387.3300 ;
      RECT 1111.2600 2381.5000 1118.7200 2394.5300 ;
      RECT 884.8600 2381.5000 1108.6600 2387.3300 ;
      RECT 870.8000 2381.5000 878.2600 2394.5300 ;
      RECT 644.4000 2381.5000 868.2000 2387.3300 ;
      RECT 630.3400 2381.5000 637.8000 2394.5300 ;
      RECT 403.9400 2381.5000 627.7400 2387.3300 ;
      RECT 389.8800 2381.5000 397.3400 2394.5300 ;
      RECT 163.3800 2381.5000 387.2800 2387.3300 ;
      RECT 3820.2800 2377.5000 3917.8400 2617.9400 ;
      RECT 3780.3800 2377.5000 3817.6800 2381.5000 ;
      RECT 3770.3800 2377.5000 3777.7800 2383.5000 ;
      RECT 3770.3800 2368.1250 3917.8400 2377.5000 ;
      RECT 3816.2800 2368.1000 3917.8400 2368.1250 ;
      RECT 3776.3800 2368.1000 3813.6800 2368.1250 ;
      RECT 3529.9200 2144.6900 3763.7800 2381.5000 ;
      RECT 3289.4600 2144.6900 3523.3200 2381.5000 ;
      RECT 3049.0000 2144.6900 3282.8600 2381.5000 ;
      RECT 2808.5400 2144.6900 3042.4000 2381.5000 ;
      RECT 2568.0800 2144.6900 2801.9400 2381.5000 ;
      RECT 2327.6200 2144.6900 2561.4800 2381.5000 ;
      RECT 2087.1600 2144.6900 2321.0200 2381.5000 ;
      RECT 1846.7000 2144.6900 2080.5600 2381.5000 ;
      RECT 1606.2400 2144.6900 1840.1000 2381.5000 ;
      RECT 1365.7800 2144.6900 1599.6400 2381.5000 ;
      RECT 1125.3200 2144.6900 1359.1800 2381.5000 ;
      RECT 884.8600 2144.6900 1118.7200 2381.5000 ;
      RECT 644.4000 2144.6900 878.2600 2381.5000 ;
      RECT 403.9400 2144.6900 637.8000 2381.5000 ;
      RECT 163.3800 2144.6900 397.3400 2381.5000 ;
      RECT 159.3800 2143.5500 160.7800 2387.3300 ;
      RECT 123.4800 2143.5500 156.7800 2388.6900 ;
      RECT 123.4800 2143.4500 150.4400 2143.5500 ;
      RECT 3816.2800 2143.2900 3817.6800 2368.1000 ;
      RECT 3780.3800 2143.2900 3813.6800 2368.1000 ;
      RECT 3780.3800 2143.1900 3807.3400 2143.2900 ;
      RECT 123.4800 2141.3500 149.7900 2143.4500 ;
      RECT 159.4800 2141.2500 160.7800 2143.5500 ;
      RECT 123.4800 2141.2500 150.4400 2141.3500 ;
      RECT 3780.3800 2141.0900 3806.6900 2143.1900 ;
      RECT 3816.3800 2140.9900 3817.6800 2143.2900 ;
      RECT 3780.3800 2140.9900 3807.3400 2141.0900 ;
      RECT 123.4800 2140.9500 156.7800 2141.2500 ;
      RECT 3780.3800 2140.7900 3813.6800 2140.9900 ;
      RECT 3776.3800 2140.7900 3777.7800 2368.1000 ;
      RECT 3784.2200 2140.6900 3813.6800 2140.7900 ;
      RECT 3529.9200 2140.2900 3753.7200 2144.6900 ;
      RECT 3525.9200 2140.2900 3527.3200 2387.3300 ;
      RECT 3289.4600 2140.2900 3513.2600 2144.6900 ;
      RECT 3285.4600 2140.2900 3286.8600 2387.3300 ;
      RECT 3049.0000 2140.2900 3272.8000 2144.6900 ;
      RECT 3045.0000 2140.2900 3046.4000 2387.3300 ;
      RECT 2808.5400 2140.2900 3032.3400 2144.6900 ;
      RECT 2804.5400 2140.2900 2805.9400 2387.3300 ;
      RECT 2568.0800 2140.2900 2791.8800 2144.6900 ;
      RECT 2564.0800 2140.2900 2565.4800 2387.3300 ;
      RECT 2327.6200 2140.2900 2551.4200 2144.6900 ;
      RECT 2323.6200 2140.2900 2325.0200 2387.3300 ;
      RECT 2087.1600 2140.2900 2310.9600 2144.6900 ;
      RECT 2083.1600 2140.2900 2084.5600 2387.3300 ;
      RECT 1846.7000 2140.2900 2070.5000 2144.6900 ;
      RECT 1842.7000 2140.2900 1844.1000 2387.3300 ;
      RECT 1606.2400 2140.2900 1830.0400 2144.6900 ;
      RECT 1602.2400 2140.2900 1603.6400 2387.3300 ;
      RECT 1365.7800 2140.2900 1589.5800 2144.6900 ;
      RECT 1361.7800 2140.2900 1363.1800 2387.3300 ;
      RECT 1125.3200 2140.2900 1349.1200 2144.6900 ;
      RECT 1121.3200 2140.2900 1122.7200 2387.3300 ;
      RECT 884.8600 2140.2900 1108.6600 2144.6900 ;
      RECT 880.8600 2140.2900 882.2600 2387.3300 ;
      RECT 644.4000 2140.2900 868.2000 2144.6900 ;
      RECT 640.4000 2140.2900 641.8000 2387.3300 ;
      RECT 403.9400 2140.2900 627.7400 2144.6900 ;
      RECT 399.9400 2140.2900 401.3400 2387.3300 ;
      RECT 163.3800 2140.2900 387.2800 2144.6900 ;
      RECT 159.3800 2140.2900 160.7800 2141.2500 ;
      RECT 3535.0800 2140.1900 3753.7200 2140.2900 ;
      RECT 3294.6200 2140.1900 3513.2600 2140.2900 ;
      RECT 3054.1600 2140.1900 3272.8000 2140.2900 ;
      RECT 2813.7000 2140.1900 3032.3400 2140.2900 ;
      RECT 2573.2400 2140.1900 2791.8800 2140.2900 ;
      RECT 2332.7800 2140.1900 2551.4200 2140.2900 ;
      RECT 2092.3200 2140.1900 2310.9600 2140.2900 ;
      RECT 1851.8600 2140.1900 2070.5000 2140.2900 ;
      RECT 1611.4000 2140.1900 1830.0400 2140.2900 ;
      RECT 1370.9400 2140.1900 1589.5800 2140.2900 ;
      RECT 1130.4800 2140.1900 1349.1200 2140.2900 ;
      RECT 890.0200 2140.1900 1108.6600 2140.2900 ;
      RECT 649.5600 2140.1900 868.2000 2140.2900 ;
      RECT 409.1000 2140.1900 627.7400 2140.2900 ;
      RECT 168.6400 2140.1900 387.2800 2140.2900 ;
      RECT 156.3100 2138.8500 156.7800 2140.9500 ;
      RECT 123.4800 2138.8500 151.7050 2140.9500 ;
      RECT 3784.8700 2138.5900 3813.6800 2140.6900 ;
      RECT 3784.2200 2138.4900 3813.6800 2138.5900 ;
      RECT 3776.3800 2138.4900 3777.6800 2140.7900 ;
      RECT 3536.4800 2137.5900 3753.7200 2140.1900 ;
      RECT 3296.0200 2137.5900 3513.2600 2140.1900 ;
      RECT 3055.5600 2137.5900 3272.8000 2140.1900 ;
      RECT 2815.1000 2137.5900 3032.3400 2140.1900 ;
      RECT 2574.6400 2137.5900 2791.8800 2140.1900 ;
      RECT 2334.1800 2137.5900 2551.4200 2140.1900 ;
      RECT 2093.7200 2137.5900 2310.9600 2140.1900 ;
      RECT 1853.2600 2137.5900 2070.5000 2140.1900 ;
      RECT 1612.8000 2137.5900 1830.0400 2140.1900 ;
      RECT 1372.3400 2137.5900 1589.5800 2140.1900 ;
      RECT 1131.8800 2137.5900 1349.1200 2140.1900 ;
      RECT 891.4200 2137.5900 1108.6600 2140.1900 ;
      RECT 650.9600 2137.5900 868.2000 2140.1900 ;
      RECT 410.5000 2137.5900 627.7400 2140.1900 ;
      RECT 170.0400 2137.5900 387.2800 2140.1900 ;
      RECT 3535.0800 2137.4900 3753.7200 2137.5900 ;
      RECT 3525.9200 2137.4900 3527.2200 2140.2900 ;
      RECT 3294.6200 2137.4900 3513.2600 2137.5900 ;
      RECT 3285.4600 2137.4900 3286.7600 2140.2900 ;
      RECT 3054.1600 2137.4900 3272.8000 2137.5900 ;
      RECT 3045.0000 2137.4900 3046.3000 2140.2900 ;
      RECT 2813.7000 2137.4900 3032.3400 2137.5900 ;
      RECT 2804.5400 2137.4900 2805.8400 2140.2900 ;
      RECT 2573.2400 2137.4900 2791.8800 2137.5900 ;
      RECT 2564.0800 2137.4900 2565.3800 2140.2900 ;
      RECT 2332.7800 2137.4900 2551.4200 2137.5900 ;
      RECT 2323.6200 2137.4900 2324.9200 2140.2900 ;
      RECT 2092.3200 2137.4900 2310.9600 2137.5900 ;
      RECT 2083.1600 2137.4900 2084.4600 2140.2900 ;
      RECT 1851.8600 2137.4900 2070.5000 2137.5900 ;
      RECT 1842.7000 2137.4900 1844.0000 2140.2900 ;
      RECT 1611.4000 2137.4900 1830.0400 2137.5900 ;
      RECT 1602.2400 2137.4900 1603.5400 2140.2900 ;
      RECT 1370.9400 2137.4900 1589.5800 2137.5900 ;
      RECT 1361.7800 2137.4900 1363.0800 2140.2900 ;
      RECT 1130.4800 2137.4900 1349.1200 2137.5900 ;
      RECT 1121.3200 2137.4900 1122.6200 2140.2900 ;
      RECT 890.0200 2137.4900 1108.6600 2137.5900 ;
      RECT 880.8600 2137.4900 882.1600 2140.2900 ;
      RECT 649.5600 2137.4900 868.2000 2137.5900 ;
      RECT 640.4000 2137.4900 641.7000 2140.2900 ;
      RECT 409.1000 2137.4900 627.7400 2137.5900 ;
      RECT 399.9400 2137.4900 401.2400 2140.2900 ;
      RECT 168.6400 2137.4900 387.2800 2137.5900 ;
      RECT 159.3800 2137.4900 160.6800 2140.2900 ;
      RECT 3776.3800 2133.6600 3777.7800 2138.4900 ;
      RECT 3770.3800 2133.6600 3773.7800 2368.1250 ;
      RECT 3816.2800 2131.6600 3817.6800 2140.9900 ;
      RECT 3780.3800 2131.6600 3813.6800 2138.4900 ;
      RECT 3756.3200 2131.6600 3763.7800 2144.6900 ;
      RECT 3529.9200 2131.6600 3753.7200 2137.4900 ;
      RECT 3515.8600 2131.6600 3523.3200 2144.6900 ;
      RECT 3289.4600 2131.6600 3513.2600 2137.4900 ;
      RECT 3275.4000 2131.6600 3282.8600 2144.6900 ;
      RECT 3049.0000 2131.6600 3272.8000 2137.4900 ;
      RECT 3034.9400 2131.6600 3042.4000 2144.6900 ;
      RECT 2808.5400 2131.6600 3032.3400 2137.4900 ;
      RECT 2794.4800 2131.6600 2801.9400 2144.6900 ;
      RECT 2568.0800 2131.6600 2791.8800 2137.4900 ;
      RECT 2554.0200 2131.6600 2561.4800 2144.6900 ;
      RECT 2327.6200 2131.6600 2551.4200 2137.4900 ;
      RECT 2313.5600 2131.6600 2321.0200 2144.6900 ;
      RECT 2087.1600 2131.6600 2310.9600 2137.4900 ;
      RECT 2073.1000 2131.6600 2080.5600 2144.6900 ;
      RECT 1846.7000 2131.6600 2070.5000 2137.4900 ;
      RECT 1832.6400 2131.6600 1840.1000 2144.6900 ;
      RECT 1606.2400 2131.6600 1830.0400 2137.4900 ;
      RECT 1592.1800 2131.6600 1599.6400 2144.6900 ;
      RECT 1365.7800 2131.6600 1589.5800 2137.4900 ;
      RECT 1351.7200 2131.6600 1359.1800 2144.6900 ;
      RECT 1125.3200 2131.6600 1349.1200 2137.4900 ;
      RECT 1111.2600 2131.6600 1118.7200 2144.6900 ;
      RECT 884.8600 2131.6600 1108.6600 2137.4900 ;
      RECT 870.8000 2131.6600 878.2600 2144.6900 ;
      RECT 644.4000 2131.6600 868.2000 2137.4900 ;
      RECT 630.3400 2131.6600 637.8000 2144.6900 ;
      RECT 403.9400 2131.6600 627.7400 2137.4900 ;
      RECT 389.8800 2131.6600 397.3400 2144.6900 ;
      RECT 163.3800 2131.6600 387.2800 2137.4900 ;
      RECT 3820.2800 2127.6600 3917.8400 2368.1000 ;
      RECT 3780.3800 2127.6600 3817.6800 2131.6600 ;
      RECT 3770.3800 2127.6600 3777.7800 2133.6600 ;
      RECT 3770.3800 2118.2600 3917.8400 2127.6600 ;
      RECT 3529.9200 1894.8500 3763.7800 2131.6600 ;
      RECT 3289.4600 1894.8500 3523.3200 2131.6600 ;
      RECT 3049.0000 1894.8500 3282.8600 2131.6600 ;
      RECT 2808.5400 1894.8500 3042.4000 2131.6600 ;
      RECT 2568.0800 1894.8500 2801.9400 2131.6600 ;
      RECT 2327.6200 1894.8500 2561.4800 2131.6600 ;
      RECT 2087.1600 1894.8500 2321.0200 2131.6600 ;
      RECT 1846.7000 1894.8500 2080.5600 2131.6600 ;
      RECT 1606.2400 1894.8500 1840.1000 2131.6600 ;
      RECT 1365.7800 1894.8500 1599.6400 2131.6600 ;
      RECT 1125.3200 1894.8500 1359.1800 2131.6600 ;
      RECT 884.8600 1894.8500 1118.7200 2131.6600 ;
      RECT 644.4000 1894.8500 878.2600 2131.6600 ;
      RECT 403.9400 1894.8500 637.8000 2131.6600 ;
      RECT 163.3800 1894.8500 397.3400 2131.6600 ;
      RECT 159.3800 1893.7100 160.7800 2137.4900 ;
      RECT 123.4800 1893.7100 156.7800 2138.8500 ;
      RECT 123.4800 1893.6100 150.4400 1893.7100 ;
      RECT 3816.2800 1893.4500 3817.6800 2118.2600 ;
      RECT 3780.3800 1893.4500 3813.6800 2118.2600 ;
      RECT 3780.3800 1893.3500 3807.3400 1893.4500 ;
      RECT 123.4800 1891.5100 149.7900 1893.6100 ;
      RECT 159.4800 1891.4100 160.7800 1893.7100 ;
      RECT 123.4800 1891.4100 150.4400 1891.5100 ;
      RECT 3780.3800 1891.2500 3806.6900 1893.3500 ;
      RECT 3816.3800 1891.1500 3817.6800 1893.4500 ;
      RECT 3780.3800 1891.1500 3807.3400 1891.2500 ;
      RECT 123.4800 1891.1100 156.7800 1891.4100 ;
      RECT 3780.3800 1890.9500 3813.6800 1891.1500 ;
      RECT 3776.3800 1890.9500 3777.7800 2118.2600 ;
      RECT 3784.2200 1890.8500 3813.6800 1890.9500 ;
      RECT 3529.9200 1890.4500 3753.7200 1894.8500 ;
      RECT 3525.9200 1890.4500 3527.3200 2137.4900 ;
      RECT 3289.4600 1890.4500 3513.2600 1894.8500 ;
      RECT 3285.4600 1890.4500 3286.8600 2137.4900 ;
      RECT 3049.0000 1890.4500 3272.8000 1894.8500 ;
      RECT 3045.0000 1890.4500 3046.4000 2137.4900 ;
      RECT 2808.5400 1890.4500 3032.3400 1894.8500 ;
      RECT 2804.5400 1890.4500 2805.9400 2137.4900 ;
      RECT 2568.0800 1890.4500 2791.8800 1894.8500 ;
      RECT 2564.0800 1890.4500 2565.4800 2137.4900 ;
      RECT 2327.6200 1890.4500 2551.4200 1894.8500 ;
      RECT 2323.6200 1890.4500 2325.0200 2137.4900 ;
      RECT 2087.1600 1890.4500 2310.9600 1894.8500 ;
      RECT 2083.1600 1890.4500 2084.5600 2137.4900 ;
      RECT 1846.7000 1890.4500 2070.5000 1894.8500 ;
      RECT 1842.7000 1890.4500 1844.1000 2137.4900 ;
      RECT 1606.2400 1890.4500 1830.0400 1894.8500 ;
      RECT 1602.2400 1890.4500 1603.6400 2137.4900 ;
      RECT 1365.7800 1890.4500 1589.5800 1894.8500 ;
      RECT 1361.7800 1890.4500 1363.1800 2137.4900 ;
      RECT 1125.3200 1890.4500 1349.1200 1894.8500 ;
      RECT 1121.3200 1890.4500 1122.7200 2137.4900 ;
      RECT 884.8600 1890.4500 1108.6600 1894.8500 ;
      RECT 880.8600 1890.4500 882.2600 2137.4900 ;
      RECT 644.4000 1890.4500 868.2000 1894.8500 ;
      RECT 640.4000 1890.4500 641.8000 2137.4900 ;
      RECT 403.9400 1890.4500 627.7400 1894.8500 ;
      RECT 399.9400 1890.4500 401.3400 2137.4900 ;
      RECT 163.3800 1890.4500 387.2800 1894.8500 ;
      RECT 159.3800 1890.4500 160.7800 1891.4100 ;
      RECT 3535.0800 1890.3500 3753.7200 1890.4500 ;
      RECT 3294.6200 1890.3500 3513.2600 1890.4500 ;
      RECT 3054.1600 1890.3500 3272.8000 1890.4500 ;
      RECT 2813.7000 1890.3500 3032.3400 1890.4500 ;
      RECT 2573.2400 1890.3500 2791.8800 1890.4500 ;
      RECT 2332.7800 1890.3500 2551.4200 1890.4500 ;
      RECT 2092.3200 1890.3500 2310.9600 1890.4500 ;
      RECT 1851.8600 1890.3500 2070.5000 1890.4500 ;
      RECT 1611.4000 1890.3500 1830.0400 1890.4500 ;
      RECT 1370.9400 1890.3500 1589.5800 1890.4500 ;
      RECT 1130.4800 1890.3500 1349.1200 1890.4500 ;
      RECT 890.0200 1890.3500 1108.6600 1890.4500 ;
      RECT 649.5600 1890.3500 868.2000 1890.4500 ;
      RECT 409.1000 1890.3500 627.7400 1890.4500 ;
      RECT 168.6400 1890.3500 387.2800 1890.4500 ;
      RECT 156.3100 1889.0100 156.7800 1891.1100 ;
      RECT 123.4800 1889.0100 151.7050 1891.1100 ;
      RECT 3784.8700 1888.7500 3813.6800 1890.8500 ;
      RECT 3784.2200 1888.6500 3813.6800 1888.7500 ;
      RECT 3776.3800 1888.6500 3777.6800 1890.9500 ;
      RECT 3536.4800 1887.7500 3753.7200 1890.3500 ;
      RECT 3296.0200 1887.7500 3513.2600 1890.3500 ;
      RECT 3055.5600 1887.7500 3272.8000 1890.3500 ;
      RECT 2815.1000 1887.7500 3032.3400 1890.3500 ;
      RECT 2574.6400 1887.7500 2791.8800 1890.3500 ;
      RECT 2334.1800 1887.7500 2551.4200 1890.3500 ;
      RECT 2093.7200 1887.7500 2310.9600 1890.3500 ;
      RECT 1853.2600 1887.7500 2070.5000 1890.3500 ;
      RECT 1612.8000 1887.7500 1830.0400 1890.3500 ;
      RECT 1372.3400 1887.7500 1589.5800 1890.3500 ;
      RECT 1131.8800 1887.7500 1349.1200 1890.3500 ;
      RECT 891.4200 1887.7500 1108.6600 1890.3500 ;
      RECT 650.9600 1887.7500 868.2000 1890.3500 ;
      RECT 410.5000 1887.7500 627.7400 1890.3500 ;
      RECT 170.0400 1887.7500 387.2800 1890.3500 ;
      RECT 3535.0800 1887.6500 3753.7200 1887.7500 ;
      RECT 3525.9200 1887.6500 3527.2200 1890.4500 ;
      RECT 3294.6200 1887.6500 3513.2600 1887.7500 ;
      RECT 3285.4600 1887.6500 3286.7600 1890.4500 ;
      RECT 3054.1600 1887.6500 3272.8000 1887.7500 ;
      RECT 3045.0000 1887.6500 3046.3000 1890.4500 ;
      RECT 2813.7000 1887.6500 3032.3400 1887.7500 ;
      RECT 2804.5400 1887.6500 2805.8400 1890.4500 ;
      RECT 2573.2400 1887.6500 2791.8800 1887.7500 ;
      RECT 2564.0800 1887.6500 2565.3800 1890.4500 ;
      RECT 2332.7800 1887.6500 2551.4200 1887.7500 ;
      RECT 2323.6200 1887.6500 2324.9200 1890.4500 ;
      RECT 2092.3200 1887.6500 2310.9600 1887.7500 ;
      RECT 2083.1600 1887.6500 2084.4600 1890.4500 ;
      RECT 1851.8600 1887.6500 2070.5000 1887.7500 ;
      RECT 1842.7000 1887.6500 1844.0000 1890.4500 ;
      RECT 1611.4000 1887.6500 1830.0400 1887.7500 ;
      RECT 1602.2400 1887.6500 1603.5400 1890.4500 ;
      RECT 1370.9400 1887.6500 1589.5800 1887.7500 ;
      RECT 1361.7800 1887.6500 1363.0800 1890.4500 ;
      RECT 1130.4800 1887.6500 1349.1200 1887.7500 ;
      RECT 1121.3200 1887.6500 1122.6200 1890.4500 ;
      RECT 890.0200 1887.6500 1108.6600 1887.7500 ;
      RECT 880.8600 1887.6500 882.1600 1890.4500 ;
      RECT 649.5600 1887.6500 868.2000 1887.7500 ;
      RECT 640.4000 1887.6500 641.7000 1890.4500 ;
      RECT 409.1000 1887.6500 627.7400 1887.7500 ;
      RECT 399.9400 1887.6500 401.2400 1890.4500 ;
      RECT 168.6400 1887.6500 387.2800 1887.7500 ;
      RECT 159.3800 1887.6500 160.6800 1890.4500 ;
      RECT 3776.3800 1883.8200 3777.7800 1888.6500 ;
      RECT 3770.3800 1883.8200 3773.7800 2118.2600 ;
      RECT 3816.2800 1881.8200 3817.6800 1891.1500 ;
      RECT 3780.3800 1881.8200 3813.6800 1888.6500 ;
      RECT 3756.3200 1881.8200 3763.7800 1894.8500 ;
      RECT 3529.9200 1881.8200 3753.7200 1887.6500 ;
      RECT 3515.8600 1881.8200 3523.3200 1894.8500 ;
      RECT 3289.4600 1881.8200 3513.2600 1887.6500 ;
      RECT 3275.4000 1881.8200 3282.8600 1894.8500 ;
      RECT 3049.0000 1881.8200 3272.8000 1887.6500 ;
      RECT 3034.9400 1881.8200 3042.4000 1894.8500 ;
      RECT 2808.5400 1881.8200 3032.3400 1887.6500 ;
      RECT 2794.4800 1881.8200 2801.9400 1894.8500 ;
      RECT 2568.0800 1881.8200 2791.8800 1887.6500 ;
      RECT 2554.0200 1881.8200 2561.4800 1894.8500 ;
      RECT 2327.6200 1881.8200 2551.4200 1887.6500 ;
      RECT 2313.5600 1881.8200 2321.0200 1894.8500 ;
      RECT 2087.1600 1881.8200 2310.9600 1887.6500 ;
      RECT 2073.1000 1881.8200 2080.5600 1894.8500 ;
      RECT 1846.7000 1881.8200 2070.5000 1887.6500 ;
      RECT 1832.6400 1881.8200 1840.1000 1894.8500 ;
      RECT 1606.2400 1881.8200 1830.0400 1887.6500 ;
      RECT 1592.1800 1881.8200 1599.6400 1894.8500 ;
      RECT 1365.7800 1881.8200 1589.5800 1887.6500 ;
      RECT 1351.7200 1881.8200 1359.1800 1894.8500 ;
      RECT 1125.3200 1881.8200 1349.1200 1887.6500 ;
      RECT 1111.2600 1881.8200 1118.7200 1894.8500 ;
      RECT 884.8600 1881.8200 1108.6600 1887.6500 ;
      RECT 870.8000 1881.8200 878.2600 1894.8500 ;
      RECT 644.4000 1881.8200 868.2000 1887.6500 ;
      RECT 630.3400 1881.8200 637.8000 1894.8500 ;
      RECT 403.9400 1881.8200 627.7400 1887.6500 ;
      RECT 389.8800 1881.8200 397.3400 1894.8500 ;
      RECT 163.3800 1881.8200 387.2800 1887.6500 ;
      RECT 3820.2800 1877.8200 3917.8400 2118.2600 ;
      RECT 3780.3800 1877.8200 3817.6800 1881.8200 ;
      RECT 3770.3800 1877.8200 3777.7800 1883.8200 ;
      RECT 3770.3800 1868.4200 3917.8400 1877.8200 ;
      RECT 3529.9200 1645.0100 3763.7800 1881.8200 ;
      RECT 3289.4600 1645.0100 3523.3200 1881.8200 ;
      RECT 3049.0000 1645.0100 3282.8600 1881.8200 ;
      RECT 2808.5400 1645.0100 3042.4000 1881.8200 ;
      RECT 2568.0800 1645.0100 2801.9400 1881.8200 ;
      RECT 2327.6200 1645.0100 2561.4800 1881.8200 ;
      RECT 2087.1600 1645.0100 2321.0200 1881.8200 ;
      RECT 1846.7000 1645.0100 2080.5600 1881.8200 ;
      RECT 1606.2400 1645.0100 1840.1000 1881.8200 ;
      RECT 1365.7800 1645.0100 1599.6400 1881.8200 ;
      RECT 1125.3200 1645.0100 1359.1800 1881.8200 ;
      RECT 884.8600 1645.0100 1118.7200 1881.8200 ;
      RECT 644.4000 1645.0100 878.2600 1881.8200 ;
      RECT 403.9400 1645.0100 637.8000 1881.8200 ;
      RECT 163.3800 1645.0100 397.3400 1881.8200 ;
      RECT 159.3800 1643.8700 160.7800 1887.6500 ;
      RECT 123.4800 1643.8700 156.7800 1889.0100 ;
      RECT 123.4800 1643.7700 150.4400 1643.8700 ;
      RECT 3816.2800 1643.6100 3817.6800 1868.4200 ;
      RECT 3780.3800 1643.6100 3813.6800 1868.4200 ;
      RECT 3780.3800 1643.5100 3807.3400 1643.6100 ;
      RECT 123.4800 1641.6700 149.7900 1643.7700 ;
      RECT 159.4800 1641.5700 160.7800 1643.8700 ;
      RECT 123.4800 1641.5700 150.4400 1641.6700 ;
      RECT 3780.3800 1641.4100 3806.6900 1643.5100 ;
      RECT 3816.3800 1641.3100 3817.6800 1643.6100 ;
      RECT 3780.3800 1641.3100 3807.3400 1641.4100 ;
      RECT 123.4800 1641.2700 156.7800 1641.5700 ;
      RECT 3780.3800 1641.1100 3813.6800 1641.3100 ;
      RECT 3776.3800 1641.1100 3777.7800 1868.4200 ;
      RECT 3784.2200 1641.0100 3813.6800 1641.1100 ;
      RECT 3529.9200 1640.6100 3753.7200 1645.0100 ;
      RECT 3525.9200 1640.6100 3527.3200 1887.6500 ;
      RECT 3289.4600 1640.6100 3513.2600 1645.0100 ;
      RECT 3285.4600 1640.6100 3286.8600 1887.6500 ;
      RECT 3049.0000 1640.6100 3272.8000 1645.0100 ;
      RECT 3045.0000 1640.6100 3046.4000 1887.6500 ;
      RECT 2808.5400 1640.6100 3032.3400 1645.0100 ;
      RECT 2804.5400 1640.6100 2805.9400 1887.6500 ;
      RECT 2568.0800 1640.6100 2791.8800 1645.0100 ;
      RECT 2564.0800 1640.6100 2565.4800 1887.6500 ;
      RECT 2327.6200 1640.6100 2551.4200 1645.0100 ;
      RECT 2323.6200 1640.6100 2325.0200 1887.6500 ;
      RECT 2087.1600 1640.6100 2310.9600 1645.0100 ;
      RECT 2083.1600 1640.6100 2084.5600 1887.6500 ;
      RECT 1846.7000 1640.6100 2070.5000 1645.0100 ;
      RECT 1842.7000 1640.6100 1844.1000 1887.6500 ;
      RECT 1606.2400 1640.6100 1830.0400 1645.0100 ;
      RECT 1602.2400 1640.6100 1603.6400 1887.6500 ;
      RECT 1365.7800 1640.6100 1589.5800 1645.0100 ;
      RECT 1361.7800 1640.6100 1363.1800 1887.6500 ;
      RECT 1125.3200 1640.6100 1349.1200 1645.0100 ;
      RECT 1121.3200 1640.6100 1122.7200 1887.6500 ;
      RECT 884.8600 1640.6100 1108.6600 1645.0100 ;
      RECT 880.8600 1640.6100 882.2600 1887.6500 ;
      RECT 644.4000 1640.6100 868.2000 1645.0100 ;
      RECT 640.4000 1640.6100 641.8000 1887.6500 ;
      RECT 403.9400 1640.6100 627.7400 1645.0100 ;
      RECT 399.9400 1640.6100 401.3400 1887.6500 ;
      RECT 163.3800 1640.6100 387.2800 1645.0100 ;
      RECT 159.3800 1640.6100 160.7800 1641.5700 ;
      RECT 3535.0800 1640.5100 3753.7200 1640.6100 ;
      RECT 3294.6200 1640.5100 3513.2600 1640.6100 ;
      RECT 3054.1600 1640.5100 3272.8000 1640.6100 ;
      RECT 2813.7000 1640.5100 3032.3400 1640.6100 ;
      RECT 2573.2400 1640.5100 2791.8800 1640.6100 ;
      RECT 2332.7800 1640.5100 2551.4200 1640.6100 ;
      RECT 2092.3200 1640.5100 2310.9600 1640.6100 ;
      RECT 1851.8600 1640.5100 2070.5000 1640.6100 ;
      RECT 1611.4000 1640.5100 1830.0400 1640.6100 ;
      RECT 1370.9400 1640.5100 1589.5800 1640.6100 ;
      RECT 1130.4800 1640.5100 1349.1200 1640.6100 ;
      RECT 890.0200 1640.5100 1108.6600 1640.6100 ;
      RECT 649.5600 1640.5100 868.2000 1640.6100 ;
      RECT 409.1000 1640.5100 627.7400 1640.6100 ;
      RECT 168.6400 1640.5100 387.2800 1640.6100 ;
      RECT 156.3100 1639.1700 156.7800 1641.2700 ;
      RECT 123.4800 1639.1700 151.7050 1641.2700 ;
      RECT 3784.8700 1638.9100 3813.6800 1641.0100 ;
      RECT 3784.2200 1638.8100 3813.6800 1638.9100 ;
      RECT 3776.3800 1638.8100 3777.6800 1641.1100 ;
      RECT 3536.4800 1637.9100 3753.7200 1640.5100 ;
      RECT 3296.0200 1637.9100 3513.2600 1640.5100 ;
      RECT 3055.5600 1637.9100 3272.8000 1640.5100 ;
      RECT 2815.1000 1637.9100 3032.3400 1640.5100 ;
      RECT 2574.6400 1637.9100 2791.8800 1640.5100 ;
      RECT 2334.1800 1637.9100 2551.4200 1640.5100 ;
      RECT 2093.7200 1637.9100 2310.9600 1640.5100 ;
      RECT 1853.2600 1637.9100 2070.5000 1640.5100 ;
      RECT 1612.8000 1637.9100 1830.0400 1640.5100 ;
      RECT 1372.3400 1637.9100 1589.5800 1640.5100 ;
      RECT 1131.8800 1637.9100 1349.1200 1640.5100 ;
      RECT 891.4200 1637.9100 1108.6600 1640.5100 ;
      RECT 650.9600 1637.9100 868.2000 1640.5100 ;
      RECT 410.5000 1637.9100 627.7400 1640.5100 ;
      RECT 170.0400 1637.9100 387.2800 1640.5100 ;
      RECT 3535.0800 1637.8100 3753.7200 1637.9100 ;
      RECT 3525.9200 1637.8100 3527.2200 1640.6100 ;
      RECT 3294.6200 1637.8100 3513.2600 1637.9100 ;
      RECT 3285.4600 1637.8100 3286.7600 1640.6100 ;
      RECT 3054.1600 1637.8100 3272.8000 1637.9100 ;
      RECT 3045.0000 1637.8100 3046.3000 1640.6100 ;
      RECT 2813.7000 1637.8100 3032.3400 1637.9100 ;
      RECT 2804.5400 1637.8100 2805.8400 1640.6100 ;
      RECT 2573.2400 1637.8100 2791.8800 1637.9100 ;
      RECT 2564.0800 1637.8100 2565.3800 1640.6100 ;
      RECT 2332.7800 1637.8100 2551.4200 1637.9100 ;
      RECT 2323.6200 1637.8100 2324.9200 1640.6100 ;
      RECT 2092.3200 1637.8100 2310.9600 1637.9100 ;
      RECT 2083.1600 1637.8100 2084.4600 1640.6100 ;
      RECT 1851.8600 1637.8100 2070.5000 1637.9100 ;
      RECT 1842.7000 1637.8100 1844.0000 1640.6100 ;
      RECT 1611.4000 1637.8100 1830.0400 1637.9100 ;
      RECT 1602.2400 1637.8100 1603.5400 1640.6100 ;
      RECT 1370.9400 1637.8100 1589.5800 1637.9100 ;
      RECT 1361.7800 1637.8100 1363.0800 1640.6100 ;
      RECT 1130.4800 1637.8100 1349.1200 1637.9100 ;
      RECT 1121.3200 1637.8100 1122.6200 1640.6100 ;
      RECT 890.0200 1637.8100 1108.6600 1637.9100 ;
      RECT 880.8600 1637.8100 882.1600 1640.6100 ;
      RECT 649.5600 1637.8100 868.2000 1637.9100 ;
      RECT 640.4000 1637.8100 641.7000 1640.6100 ;
      RECT 409.1000 1637.8100 627.7400 1637.9100 ;
      RECT 399.9400 1637.8100 401.2400 1640.6100 ;
      RECT 168.6400 1637.8100 387.2800 1637.9100 ;
      RECT 159.3800 1637.8100 160.6800 1640.6100 ;
      RECT 3776.3800 1633.9800 3777.7800 1638.8100 ;
      RECT 3770.3800 1633.9800 3773.7800 1868.4200 ;
      RECT 3816.2800 1631.9800 3817.6800 1641.3100 ;
      RECT 3780.3800 1631.9800 3813.6800 1638.8100 ;
      RECT 3756.3200 1631.9800 3763.7800 1645.0100 ;
      RECT 3529.9200 1631.9800 3753.7200 1637.8100 ;
      RECT 3515.8600 1631.9800 3523.3200 1645.0100 ;
      RECT 3289.4600 1631.9800 3513.2600 1637.8100 ;
      RECT 3275.4000 1631.9800 3282.8600 1645.0100 ;
      RECT 3049.0000 1631.9800 3272.8000 1637.8100 ;
      RECT 3034.9400 1631.9800 3042.4000 1645.0100 ;
      RECT 2808.5400 1631.9800 3032.3400 1637.8100 ;
      RECT 2794.4800 1631.9800 2801.9400 1645.0100 ;
      RECT 2568.0800 1631.9800 2791.8800 1637.8100 ;
      RECT 2554.0200 1631.9800 2561.4800 1645.0100 ;
      RECT 2327.6200 1631.9800 2551.4200 1637.8100 ;
      RECT 2313.5600 1631.9800 2321.0200 1645.0100 ;
      RECT 2087.1600 1631.9800 2310.9600 1637.8100 ;
      RECT 2073.1000 1631.9800 2080.5600 1645.0100 ;
      RECT 1846.7000 1631.9800 2070.5000 1637.8100 ;
      RECT 1832.6400 1631.9800 1840.1000 1645.0100 ;
      RECT 1606.2400 1631.9800 1830.0400 1637.8100 ;
      RECT 1592.1800 1631.9800 1599.6400 1645.0100 ;
      RECT 1365.7800 1631.9800 1589.5800 1637.8100 ;
      RECT 1351.7200 1631.9800 1359.1800 1645.0100 ;
      RECT 1125.3200 1631.9800 1349.1200 1637.8100 ;
      RECT 1111.2600 1631.9800 1118.7200 1645.0100 ;
      RECT 884.8600 1631.9800 1108.6600 1637.8100 ;
      RECT 870.8000 1631.9800 878.2600 1645.0100 ;
      RECT 644.4000 1631.9800 868.2000 1637.8100 ;
      RECT 630.3400 1631.9800 637.8000 1645.0100 ;
      RECT 403.9400 1631.9800 627.7400 1637.8100 ;
      RECT 389.8800 1631.9800 397.3400 1645.0100 ;
      RECT 163.3800 1631.9800 387.2800 1637.8100 ;
      RECT 3820.2800 1627.9800 3917.8400 1868.4200 ;
      RECT 3780.3800 1627.9800 3817.6800 1631.9800 ;
      RECT 3770.3800 1627.9800 3777.7800 1633.9800 ;
      RECT 3770.3800 1618.5800 3917.8400 1627.9800 ;
      RECT 3529.9200 1395.1700 3763.7800 1631.9800 ;
      RECT 3289.4600 1395.1700 3523.3200 1631.9800 ;
      RECT 3049.0000 1395.1700 3282.8600 1631.9800 ;
      RECT 2808.5400 1395.1700 3042.4000 1631.9800 ;
      RECT 2568.0800 1395.1700 2801.9400 1631.9800 ;
      RECT 2327.6200 1395.1700 2561.4800 1631.9800 ;
      RECT 2087.1600 1395.1700 2321.0200 1631.9800 ;
      RECT 1846.7000 1395.1700 2080.5600 1631.9800 ;
      RECT 1606.2400 1395.1700 1840.1000 1631.9800 ;
      RECT 1365.7800 1395.1700 1599.6400 1631.9800 ;
      RECT 1125.3200 1395.1700 1359.1800 1631.9800 ;
      RECT 884.8600 1395.1700 1118.7200 1631.9800 ;
      RECT 644.4000 1395.1700 878.2600 1631.9800 ;
      RECT 403.9400 1395.1700 637.8000 1631.9800 ;
      RECT 163.3800 1395.1700 397.3400 1631.9800 ;
      RECT 159.3800 1394.0300 160.7800 1637.8100 ;
      RECT 123.4800 1394.0300 156.7800 1639.1700 ;
      RECT 123.4800 1393.9300 150.4400 1394.0300 ;
      RECT 3816.2800 1393.7700 3817.6800 1618.5800 ;
      RECT 3780.3800 1393.7700 3813.6800 1618.5800 ;
      RECT 3780.3800 1393.6700 3807.3400 1393.7700 ;
      RECT 123.4800 1391.8300 149.7900 1393.9300 ;
      RECT 159.4800 1391.7300 160.7800 1394.0300 ;
      RECT 123.4800 1391.7300 150.4400 1391.8300 ;
      RECT 3780.3800 1391.5700 3806.6900 1393.6700 ;
      RECT 3816.3800 1391.4700 3817.6800 1393.7700 ;
      RECT 3780.3800 1391.4700 3807.3400 1391.5700 ;
      RECT 123.4800 1391.4300 156.7800 1391.7300 ;
      RECT 3780.3800 1391.2700 3813.6800 1391.4700 ;
      RECT 3776.3800 1391.2700 3777.7800 1618.5800 ;
      RECT 3784.2200 1391.1700 3813.6800 1391.2700 ;
      RECT 3529.9200 1390.7700 3753.7200 1395.1700 ;
      RECT 3525.9200 1390.7700 3527.3200 1637.8100 ;
      RECT 3289.4600 1390.7700 3513.2600 1395.1700 ;
      RECT 3285.4600 1390.7700 3286.8600 1637.8100 ;
      RECT 3049.0000 1390.7700 3272.8000 1395.1700 ;
      RECT 3045.0000 1390.7700 3046.4000 1637.8100 ;
      RECT 2808.5400 1390.7700 3032.3400 1395.1700 ;
      RECT 2804.5400 1390.7700 2805.9400 1637.8100 ;
      RECT 2568.0800 1390.7700 2791.8800 1395.1700 ;
      RECT 2564.0800 1390.7700 2565.4800 1637.8100 ;
      RECT 2327.6200 1390.7700 2551.4200 1395.1700 ;
      RECT 2323.6200 1390.7700 2325.0200 1637.8100 ;
      RECT 2087.1600 1390.7700 2310.9600 1395.1700 ;
      RECT 2083.1600 1390.7700 2084.5600 1637.8100 ;
      RECT 1846.7000 1390.7700 2070.5000 1395.1700 ;
      RECT 1842.7000 1390.7700 1844.1000 1637.8100 ;
      RECT 1606.2400 1390.7700 1830.0400 1395.1700 ;
      RECT 1602.2400 1390.7700 1603.6400 1637.8100 ;
      RECT 1365.7800 1390.7700 1589.5800 1395.1700 ;
      RECT 1361.7800 1390.7700 1363.1800 1637.8100 ;
      RECT 1125.3200 1390.7700 1349.1200 1395.1700 ;
      RECT 1121.3200 1390.7700 1122.7200 1637.8100 ;
      RECT 884.8600 1390.7700 1108.6600 1395.1700 ;
      RECT 880.8600 1390.7700 882.2600 1637.8100 ;
      RECT 644.4000 1390.7700 868.2000 1395.1700 ;
      RECT 640.4000 1390.7700 641.8000 1637.8100 ;
      RECT 403.9400 1390.7700 627.7400 1395.1700 ;
      RECT 399.9400 1390.7700 401.3400 1637.8100 ;
      RECT 163.3800 1390.7700 387.2800 1395.1700 ;
      RECT 159.3800 1390.7700 160.7800 1391.7300 ;
      RECT 3535.0800 1390.6700 3753.7200 1390.7700 ;
      RECT 3294.6200 1390.6700 3513.2600 1390.7700 ;
      RECT 3054.1600 1390.6700 3272.8000 1390.7700 ;
      RECT 2813.7000 1390.6700 3032.3400 1390.7700 ;
      RECT 2573.2400 1390.6700 2791.8800 1390.7700 ;
      RECT 2332.7800 1390.6700 2551.4200 1390.7700 ;
      RECT 2092.3200 1390.6700 2310.9600 1390.7700 ;
      RECT 1851.8600 1390.6700 2070.5000 1390.7700 ;
      RECT 1611.4000 1390.6700 1830.0400 1390.7700 ;
      RECT 1370.9400 1390.6700 1589.5800 1390.7700 ;
      RECT 1130.4800 1390.6700 1349.1200 1390.7700 ;
      RECT 890.0200 1390.6700 1108.6600 1390.7700 ;
      RECT 649.5600 1390.6700 868.2000 1390.7700 ;
      RECT 409.1000 1390.6700 627.7400 1390.7700 ;
      RECT 168.6400 1390.6700 387.2800 1390.7700 ;
      RECT 156.3100 1389.3300 156.7800 1391.4300 ;
      RECT 123.4800 1389.3300 151.7050 1391.4300 ;
      RECT 3784.8700 1389.0700 3813.6800 1391.1700 ;
      RECT 3784.2200 1388.9700 3813.6800 1389.0700 ;
      RECT 3776.3800 1388.9700 3777.6800 1391.2700 ;
      RECT 3536.4800 1388.0700 3753.7200 1390.6700 ;
      RECT 3296.0200 1388.0700 3513.2600 1390.6700 ;
      RECT 3055.5600 1388.0700 3272.8000 1390.6700 ;
      RECT 2815.1000 1388.0700 3032.3400 1390.6700 ;
      RECT 2574.6400 1388.0700 2791.8800 1390.6700 ;
      RECT 2334.1800 1388.0700 2551.4200 1390.6700 ;
      RECT 2093.7200 1388.0700 2310.9600 1390.6700 ;
      RECT 1853.2600 1388.0700 2070.5000 1390.6700 ;
      RECT 1612.8000 1388.0700 1830.0400 1390.6700 ;
      RECT 1372.3400 1388.0700 1589.5800 1390.6700 ;
      RECT 1131.8800 1388.0700 1349.1200 1390.6700 ;
      RECT 891.4200 1388.0700 1108.6600 1390.6700 ;
      RECT 650.9600 1388.0700 868.2000 1390.6700 ;
      RECT 410.5000 1388.0700 627.7400 1390.6700 ;
      RECT 170.0400 1388.0700 387.2800 1390.6700 ;
      RECT 3535.0800 1387.9700 3753.7200 1388.0700 ;
      RECT 3525.9200 1387.9700 3527.2200 1390.7700 ;
      RECT 3294.6200 1387.9700 3513.2600 1388.0700 ;
      RECT 3285.4600 1387.9700 3286.7600 1390.7700 ;
      RECT 3054.1600 1387.9700 3272.8000 1388.0700 ;
      RECT 3045.0000 1387.9700 3046.3000 1390.7700 ;
      RECT 2813.7000 1387.9700 3032.3400 1388.0700 ;
      RECT 2804.5400 1387.9700 2805.8400 1390.7700 ;
      RECT 2573.2400 1387.9700 2791.8800 1388.0700 ;
      RECT 2564.0800 1387.9700 2565.3800 1390.7700 ;
      RECT 2332.7800 1387.9700 2551.4200 1388.0700 ;
      RECT 2323.6200 1387.9700 2324.9200 1390.7700 ;
      RECT 2092.3200 1387.9700 2310.9600 1388.0700 ;
      RECT 2083.1600 1387.9700 2084.4600 1390.7700 ;
      RECT 1851.8600 1387.9700 2070.5000 1388.0700 ;
      RECT 1842.7000 1387.9700 1844.0000 1390.7700 ;
      RECT 1611.4000 1387.9700 1830.0400 1388.0700 ;
      RECT 1602.2400 1387.9700 1603.5400 1390.7700 ;
      RECT 1370.9400 1387.9700 1589.5800 1388.0700 ;
      RECT 1361.7800 1387.9700 1363.0800 1390.7700 ;
      RECT 1130.4800 1387.9700 1349.1200 1388.0700 ;
      RECT 1121.3200 1387.9700 1122.6200 1390.7700 ;
      RECT 890.0200 1387.9700 1108.6600 1388.0700 ;
      RECT 880.8600 1387.9700 882.1600 1390.7700 ;
      RECT 649.5600 1387.9700 868.2000 1388.0700 ;
      RECT 640.4000 1387.9700 641.7000 1390.7700 ;
      RECT 409.1000 1387.9700 627.7400 1388.0700 ;
      RECT 399.9400 1387.9700 401.2400 1390.7700 ;
      RECT 168.6400 1387.9700 387.2800 1388.0700 ;
      RECT 159.3800 1387.9700 160.6800 1390.7700 ;
      RECT 3776.3800 1384.1400 3777.7800 1388.9700 ;
      RECT 3770.3800 1384.1400 3773.7800 1618.5800 ;
      RECT 3816.2800 1382.1400 3817.6800 1391.4700 ;
      RECT 3780.3800 1382.1400 3813.6800 1388.9700 ;
      RECT 3756.3200 1382.1400 3763.7800 1395.1700 ;
      RECT 3529.9200 1382.1400 3753.7200 1387.9700 ;
      RECT 3515.8600 1382.1400 3523.3200 1395.1700 ;
      RECT 3289.4600 1382.1400 3513.2600 1387.9700 ;
      RECT 3275.4000 1382.1400 3282.8600 1395.1700 ;
      RECT 3049.0000 1382.1400 3272.8000 1387.9700 ;
      RECT 3034.9400 1382.1400 3042.4000 1395.1700 ;
      RECT 2808.5400 1382.1400 3032.3400 1387.9700 ;
      RECT 2794.4800 1382.1400 2801.9400 1395.1700 ;
      RECT 2568.0800 1382.1400 2791.8800 1387.9700 ;
      RECT 2554.0200 1382.1400 2561.4800 1395.1700 ;
      RECT 2327.6200 1382.1400 2551.4200 1387.9700 ;
      RECT 2313.5600 1382.1400 2321.0200 1395.1700 ;
      RECT 2087.1600 1382.1400 2310.9600 1387.9700 ;
      RECT 2073.1000 1382.1400 2080.5600 1395.1700 ;
      RECT 1846.7000 1382.1400 2070.5000 1387.9700 ;
      RECT 1832.6400 1382.1400 1840.1000 1395.1700 ;
      RECT 1606.2400 1382.1400 1830.0400 1387.9700 ;
      RECT 1592.1800 1382.1400 1599.6400 1395.1700 ;
      RECT 1365.7800 1382.1400 1589.5800 1387.9700 ;
      RECT 1351.7200 1382.1400 1359.1800 1395.1700 ;
      RECT 1125.3200 1382.1400 1349.1200 1387.9700 ;
      RECT 1111.2600 1382.1400 1118.7200 1395.1700 ;
      RECT 884.8600 1382.1400 1108.6600 1387.9700 ;
      RECT 870.8000 1382.1400 878.2600 1395.1700 ;
      RECT 644.4000 1382.1400 868.2000 1387.9700 ;
      RECT 630.3400 1382.1400 637.8000 1395.1700 ;
      RECT 403.9400 1382.1400 627.7400 1387.9700 ;
      RECT 389.8800 1382.1400 397.3400 1395.1700 ;
      RECT 163.3800 1382.1400 387.2800 1387.9700 ;
      RECT 3820.2800 1378.1400 3917.8400 1618.5800 ;
      RECT 3780.3800 1378.1400 3817.6800 1382.1400 ;
      RECT 3770.3800 1378.1400 3777.7800 1384.1400 ;
      RECT 3770.3800 1368.7400 3917.8400 1378.1400 ;
      RECT 3529.9200 1145.3300 3763.7800 1382.1400 ;
      RECT 3289.4600 1145.3300 3523.3200 1382.1400 ;
      RECT 3049.0000 1145.3300 3282.8600 1382.1400 ;
      RECT 2808.5400 1145.3300 3042.4000 1382.1400 ;
      RECT 2568.0800 1145.3300 2801.9400 1382.1400 ;
      RECT 2327.6200 1145.3300 2561.4800 1382.1400 ;
      RECT 2087.1600 1145.3300 2321.0200 1382.1400 ;
      RECT 1846.7000 1145.3300 2080.5600 1382.1400 ;
      RECT 1606.2400 1145.3300 1840.1000 1382.1400 ;
      RECT 1365.7800 1145.3300 1599.6400 1382.1400 ;
      RECT 1125.3200 1145.3300 1359.1800 1382.1400 ;
      RECT 884.8600 1145.3300 1118.7200 1382.1400 ;
      RECT 644.4000 1145.3300 878.2600 1382.1400 ;
      RECT 403.9400 1145.3300 637.8000 1382.1400 ;
      RECT 163.3800 1145.3300 397.3400 1382.1400 ;
      RECT 159.3800 1144.1900 160.7800 1387.9700 ;
      RECT 123.4800 1144.1900 156.7800 1389.3300 ;
      RECT 123.4800 1144.0900 150.4400 1144.1900 ;
      RECT 3816.2800 1143.9300 3817.6800 1368.7400 ;
      RECT 3780.3800 1143.9300 3813.6800 1368.7400 ;
      RECT 3780.3800 1143.8300 3807.3400 1143.9300 ;
      RECT 123.4800 1141.9900 149.7900 1144.0900 ;
      RECT 159.4800 1141.8900 160.7800 1144.1900 ;
      RECT 123.4800 1141.8900 150.4400 1141.9900 ;
      RECT 3780.3800 1141.7300 3806.6900 1143.8300 ;
      RECT 3816.3800 1141.6300 3817.6800 1143.9300 ;
      RECT 3780.3800 1141.6300 3807.3400 1141.7300 ;
      RECT 123.4800 1141.5900 156.7800 1141.8900 ;
      RECT 3780.3800 1141.4300 3813.6800 1141.6300 ;
      RECT 3776.3800 1141.4300 3777.7800 1368.7400 ;
      RECT 3784.2200 1141.3300 3813.6800 1141.4300 ;
      RECT 3529.9200 1140.9300 3753.7200 1145.3300 ;
      RECT 3525.9200 1140.9300 3527.3200 1387.9700 ;
      RECT 3289.4600 1140.9300 3513.2600 1145.3300 ;
      RECT 3285.4600 1140.9300 3286.8600 1387.9700 ;
      RECT 3049.0000 1140.9300 3272.8000 1145.3300 ;
      RECT 3045.0000 1140.9300 3046.4000 1387.9700 ;
      RECT 2808.5400 1140.9300 3032.3400 1145.3300 ;
      RECT 2804.5400 1140.9300 2805.9400 1387.9700 ;
      RECT 2568.0800 1140.9300 2791.8800 1145.3300 ;
      RECT 2564.0800 1140.9300 2565.4800 1387.9700 ;
      RECT 2327.6200 1140.9300 2551.4200 1145.3300 ;
      RECT 2323.6200 1140.9300 2325.0200 1387.9700 ;
      RECT 2087.1600 1140.9300 2310.9600 1145.3300 ;
      RECT 2083.1600 1140.9300 2084.5600 1387.9700 ;
      RECT 1846.7000 1140.9300 2070.5000 1145.3300 ;
      RECT 1842.7000 1140.9300 1844.1000 1387.9700 ;
      RECT 1606.2400 1140.9300 1830.0400 1145.3300 ;
      RECT 1602.2400 1140.9300 1603.6400 1387.9700 ;
      RECT 1365.7800 1140.9300 1589.5800 1145.3300 ;
      RECT 1361.7800 1140.9300 1363.1800 1387.9700 ;
      RECT 1125.3200 1140.9300 1349.1200 1145.3300 ;
      RECT 1121.3200 1140.9300 1122.7200 1387.9700 ;
      RECT 884.8600 1140.9300 1108.6600 1145.3300 ;
      RECT 880.8600 1140.9300 882.2600 1387.9700 ;
      RECT 644.4000 1140.9300 868.2000 1145.3300 ;
      RECT 640.4000 1140.9300 641.8000 1387.9700 ;
      RECT 403.9400 1140.9300 627.7400 1145.3300 ;
      RECT 399.9400 1140.9300 401.3400 1387.9700 ;
      RECT 163.3800 1140.9300 387.2800 1145.3300 ;
      RECT 159.3800 1140.9300 160.7800 1141.8900 ;
      RECT 3535.0800 1140.8300 3753.7200 1140.9300 ;
      RECT 3294.6200 1140.8300 3513.2600 1140.9300 ;
      RECT 3054.1600 1140.8300 3272.8000 1140.9300 ;
      RECT 2813.7000 1140.8300 3032.3400 1140.9300 ;
      RECT 2573.2400 1140.8300 2791.8800 1140.9300 ;
      RECT 2332.7800 1140.8300 2551.4200 1140.9300 ;
      RECT 2092.3200 1140.8300 2310.9600 1140.9300 ;
      RECT 1851.8600 1140.8300 2070.5000 1140.9300 ;
      RECT 1611.4000 1140.8300 1830.0400 1140.9300 ;
      RECT 1370.9400 1140.8300 1589.5800 1140.9300 ;
      RECT 1130.4800 1140.8300 1349.1200 1140.9300 ;
      RECT 890.0200 1140.8300 1108.6600 1140.9300 ;
      RECT 649.5600 1140.8300 868.2000 1140.9300 ;
      RECT 409.1000 1140.8300 627.7400 1140.9300 ;
      RECT 168.6400 1140.8300 387.2800 1140.9300 ;
      RECT 156.3100 1139.4900 156.7800 1141.5900 ;
      RECT 123.4800 1139.4900 151.7050 1141.5900 ;
      RECT 3784.8700 1139.2300 3813.6800 1141.3300 ;
      RECT 3784.2200 1139.1300 3813.6800 1139.2300 ;
      RECT 3776.3800 1139.1300 3777.6800 1141.4300 ;
      RECT 3536.4800 1138.2300 3753.7200 1140.8300 ;
      RECT 3296.0200 1138.2300 3513.2600 1140.8300 ;
      RECT 3055.5600 1138.2300 3272.8000 1140.8300 ;
      RECT 2815.1000 1138.2300 3032.3400 1140.8300 ;
      RECT 2574.6400 1138.2300 2791.8800 1140.8300 ;
      RECT 2334.1800 1138.2300 2551.4200 1140.8300 ;
      RECT 2093.7200 1138.2300 2310.9600 1140.8300 ;
      RECT 1853.2600 1138.2300 2070.5000 1140.8300 ;
      RECT 1612.8000 1138.2300 1830.0400 1140.8300 ;
      RECT 1372.3400 1138.2300 1589.5800 1140.8300 ;
      RECT 1131.8800 1138.2300 1349.1200 1140.8300 ;
      RECT 891.4200 1138.2300 1108.6600 1140.8300 ;
      RECT 650.9600 1138.2300 868.2000 1140.8300 ;
      RECT 410.5000 1138.2300 627.7400 1140.8300 ;
      RECT 170.0400 1138.2300 387.2800 1140.8300 ;
      RECT 3535.0800 1138.1300 3753.7200 1138.2300 ;
      RECT 3525.9200 1138.1300 3527.2200 1140.9300 ;
      RECT 3294.6200 1138.1300 3513.2600 1138.2300 ;
      RECT 3285.4600 1138.1300 3286.7600 1140.9300 ;
      RECT 3054.1600 1138.1300 3272.8000 1138.2300 ;
      RECT 3045.0000 1138.1300 3046.3000 1140.9300 ;
      RECT 2813.7000 1138.1300 3032.3400 1138.2300 ;
      RECT 2804.5400 1138.1300 2805.8400 1140.9300 ;
      RECT 2573.2400 1138.1300 2791.8800 1138.2300 ;
      RECT 2564.0800 1138.1300 2565.3800 1140.9300 ;
      RECT 2332.7800 1138.1300 2551.4200 1138.2300 ;
      RECT 2323.6200 1138.1300 2324.9200 1140.9300 ;
      RECT 2092.3200 1138.1300 2310.9600 1138.2300 ;
      RECT 2083.1600 1138.1300 2084.4600 1140.9300 ;
      RECT 1851.8600 1138.1300 2070.5000 1138.2300 ;
      RECT 1842.7000 1138.1300 1844.0000 1140.9300 ;
      RECT 1611.4000 1138.1300 1830.0400 1138.2300 ;
      RECT 1602.2400 1138.1300 1603.5400 1140.9300 ;
      RECT 1370.9400 1138.1300 1589.5800 1138.2300 ;
      RECT 1361.7800 1138.1300 1363.0800 1140.9300 ;
      RECT 1130.4800 1138.1300 1349.1200 1138.2300 ;
      RECT 1121.3200 1138.1300 1122.6200 1140.9300 ;
      RECT 890.0200 1138.1300 1108.6600 1138.2300 ;
      RECT 880.8600 1138.1300 882.1600 1140.9300 ;
      RECT 649.5600 1138.1300 868.2000 1138.2300 ;
      RECT 640.4000 1138.1300 641.7000 1140.9300 ;
      RECT 409.1000 1138.1300 627.7400 1138.2300 ;
      RECT 399.9400 1138.1300 401.2400 1140.9300 ;
      RECT 168.6400 1138.1300 387.2800 1138.2300 ;
      RECT 159.3800 1138.1300 160.6800 1140.9300 ;
      RECT 3776.3800 1134.3000 3777.7800 1139.1300 ;
      RECT 3770.3800 1134.3000 3773.7800 1368.7400 ;
      RECT 3816.2800 1132.3000 3817.6800 1141.6300 ;
      RECT 3780.3800 1132.3000 3813.6800 1139.1300 ;
      RECT 3756.3200 1132.3000 3763.7800 1145.3300 ;
      RECT 3529.9200 1132.3000 3753.7200 1138.1300 ;
      RECT 3515.8600 1132.3000 3523.3200 1145.3300 ;
      RECT 3289.4600 1132.3000 3513.2600 1138.1300 ;
      RECT 3275.4000 1132.3000 3282.8600 1145.3300 ;
      RECT 3049.0000 1132.3000 3272.8000 1138.1300 ;
      RECT 3034.9400 1132.3000 3042.4000 1145.3300 ;
      RECT 2808.5400 1132.3000 3032.3400 1138.1300 ;
      RECT 2794.4800 1132.3000 2801.9400 1145.3300 ;
      RECT 2568.0800 1132.3000 2791.8800 1138.1300 ;
      RECT 2554.0200 1132.3000 2561.4800 1145.3300 ;
      RECT 2327.6200 1132.3000 2551.4200 1138.1300 ;
      RECT 2313.5600 1132.3000 2321.0200 1145.3300 ;
      RECT 2087.1600 1132.3000 2310.9600 1138.1300 ;
      RECT 2073.1000 1132.3000 2080.5600 1145.3300 ;
      RECT 1846.7000 1132.3000 2070.5000 1138.1300 ;
      RECT 1832.6400 1132.3000 1840.1000 1145.3300 ;
      RECT 1606.2400 1132.3000 1830.0400 1138.1300 ;
      RECT 1592.1800 1132.3000 1599.6400 1145.3300 ;
      RECT 1365.7800 1132.3000 1589.5800 1138.1300 ;
      RECT 1351.7200 1132.3000 1359.1800 1145.3300 ;
      RECT 1125.3200 1132.3000 1349.1200 1138.1300 ;
      RECT 1111.2600 1132.3000 1118.7200 1145.3300 ;
      RECT 884.8600 1132.3000 1108.6600 1138.1300 ;
      RECT 870.8000 1132.3000 878.2600 1145.3300 ;
      RECT 644.4000 1132.3000 868.2000 1138.1300 ;
      RECT 630.3400 1132.3000 637.8000 1145.3300 ;
      RECT 403.9400 1132.3000 627.7400 1138.1300 ;
      RECT 389.8800 1132.3000 397.3400 1145.3300 ;
      RECT 163.3800 1132.3000 387.2800 1138.1300 ;
      RECT 3820.2800 1128.3000 3917.8400 1368.7400 ;
      RECT 3780.3800 1128.3000 3817.6800 1132.3000 ;
      RECT 3770.3800 1128.3000 3777.7800 1134.3000 ;
      RECT 3770.3800 1118.9000 3917.8400 1128.3000 ;
      RECT 3529.9200 895.4900 3763.7800 1132.3000 ;
      RECT 3289.4600 895.4900 3523.3200 1132.3000 ;
      RECT 3049.0000 895.4900 3282.8600 1132.3000 ;
      RECT 2808.5400 895.4900 3042.4000 1132.3000 ;
      RECT 2568.0800 895.4900 2801.9400 1132.3000 ;
      RECT 2327.6200 895.4900 2561.4800 1132.3000 ;
      RECT 2087.1600 895.4900 2321.0200 1132.3000 ;
      RECT 1846.7000 895.4900 2080.5600 1132.3000 ;
      RECT 1606.2400 895.4900 1840.1000 1132.3000 ;
      RECT 1365.7800 895.4900 1599.6400 1132.3000 ;
      RECT 1125.3200 895.4900 1359.1800 1132.3000 ;
      RECT 884.8600 895.4900 1118.7200 1132.3000 ;
      RECT 644.4000 895.4900 878.2600 1132.3000 ;
      RECT 403.9400 895.4900 637.8000 1132.3000 ;
      RECT 163.3800 895.4900 397.3400 1132.3000 ;
      RECT 159.3800 894.3500 160.7800 1138.1300 ;
      RECT 123.4800 894.3500 156.7800 1139.4900 ;
      RECT 123.4800 894.2500 150.4400 894.3500 ;
      RECT 3816.2800 894.0900 3817.6800 1118.9000 ;
      RECT 3780.3800 894.0900 3813.6800 1118.9000 ;
      RECT 3780.3800 893.9900 3807.3400 894.0900 ;
      RECT 123.4800 892.1500 149.7900 894.2500 ;
      RECT 159.4800 892.0500 160.7800 894.3500 ;
      RECT 123.4800 892.0500 150.4400 892.1500 ;
      RECT 3780.3800 891.8900 3806.6900 893.9900 ;
      RECT 3816.3800 891.7900 3817.6800 894.0900 ;
      RECT 3780.3800 891.7900 3807.3400 891.8900 ;
      RECT 123.4800 891.7500 156.7800 892.0500 ;
      RECT 3780.3800 891.5900 3813.6800 891.7900 ;
      RECT 3776.3800 891.5900 3777.7800 1118.9000 ;
      RECT 3784.2200 891.4900 3813.6800 891.5900 ;
      RECT 3529.9200 891.0900 3753.7200 895.4900 ;
      RECT 3525.9200 891.0900 3527.3200 1138.1300 ;
      RECT 3289.4600 891.0900 3513.2600 895.4900 ;
      RECT 3285.4600 891.0900 3286.8600 1138.1300 ;
      RECT 3049.0000 891.0900 3272.8000 895.4900 ;
      RECT 3045.0000 891.0900 3046.4000 1138.1300 ;
      RECT 2808.5400 891.0900 3032.3400 895.4900 ;
      RECT 2804.5400 891.0900 2805.9400 1138.1300 ;
      RECT 2568.0800 891.0900 2791.8800 895.4900 ;
      RECT 2564.0800 891.0900 2565.4800 1138.1300 ;
      RECT 2327.6200 891.0900 2551.4200 895.4900 ;
      RECT 2323.6200 891.0900 2325.0200 1138.1300 ;
      RECT 2087.1600 891.0900 2310.9600 895.4900 ;
      RECT 2083.1600 891.0900 2084.5600 1138.1300 ;
      RECT 1846.7000 891.0900 2070.5000 895.4900 ;
      RECT 1842.7000 891.0900 1844.1000 1138.1300 ;
      RECT 1606.2400 891.0900 1830.0400 895.4900 ;
      RECT 1602.2400 891.0900 1603.6400 1138.1300 ;
      RECT 1365.7800 891.0900 1589.5800 895.4900 ;
      RECT 1361.7800 891.0900 1363.1800 1138.1300 ;
      RECT 1125.3200 891.0900 1349.1200 895.4900 ;
      RECT 1121.3200 891.0900 1122.7200 1138.1300 ;
      RECT 884.8600 891.0900 1108.6600 895.4900 ;
      RECT 880.8600 891.0900 882.2600 1138.1300 ;
      RECT 644.4000 891.0900 868.2000 895.4900 ;
      RECT 640.4000 891.0900 641.8000 1138.1300 ;
      RECT 403.9400 891.0900 627.7400 895.4900 ;
      RECT 399.9400 891.0900 401.3400 1138.1300 ;
      RECT 163.3800 891.0900 387.2800 895.4900 ;
      RECT 159.3800 891.0900 160.7800 892.0500 ;
      RECT 3535.0800 890.9900 3753.7200 891.0900 ;
      RECT 3294.6200 890.9900 3513.2600 891.0900 ;
      RECT 3054.1600 890.9900 3272.8000 891.0900 ;
      RECT 2813.7000 890.9900 3032.3400 891.0900 ;
      RECT 2573.2400 890.9900 2791.8800 891.0900 ;
      RECT 2332.7800 890.9900 2551.4200 891.0900 ;
      RECT 2092.3200 890.9900 2310.9600 891.0900 ;
      RECT 1851.8600 890.9900 2070.5000 891.0900 ;
      RECT 1611.4000 890.9900 1830.0400 891.0900 ;
      RECT 1370.9400 890.9900 1589.5800 891.0900 ;
      RECT 1130.4800 890.9900 1349.1200 891.0900 ;
      RECT 890.0200 890.9900 1108.6600 891.0900 ;
      RECT 649.5600 890.9900 868.2000 891.0900 ;
      RECT 409.1000 890.9900 627.7400 891.0900 ;
      RECT 168.6400 890.9900 387.2800 891.0900 ;
      RECT 156.3100 889.6500 156.7800 891.7500 ;
      RECT 123.4800 889.6500 151.7050 891.7500 ;
      RECT 3784.8700 889.3900 3813.6800 891.4900 ;
      RECT 3784.2200 889.2900 3813.6800 889.3900 ;
      RECT 3776.3800 889.2900 3777.6800 891.5900 ;
      RECT 3536.4800 888.3900 3753.7200 890.9900 ;
      RECT 3296.0200 888.3900 3513.2600 890.9900 ;
      RECT 3055.5600 888.3900 3272.8000 890.9900 ;
      RECT 2815.1000 888.3900 3032.3400 890.9900 ;
      RECT 2574.6400 888.3900 2791.8800 890.9900 ;
      RECT 2334.1800 888.3900 2551.4200 890.9900 ;
      RECT 2093.7200 888.3900 2310.9600 890.9900 ;
      RECT 1853.2600 888.3900 2070.5000 890.9900 ;
      RECT 1612.8000 888.3900 1830.0400 890.9900 ;
      RECT 1372.3400 888.3900 1589.5800 890.9900 ;
      RECT 1131.8800 888.3900 1349.1200 890.9900 ;
      RECT 891.4200 888.3900 1108.6600 890.9900 ;
      RECT 650.9600 888.3900 868.2000 890.9900 ;
      RECT 410.5000 888.3900 627.7400 890.9900 ;
      RECT 170.0400 888.3900 387.2800 890.9900 ;
      RECT 3535.0800 888.2900 3753.7200 888.3900 ;
      RECT 3525.9200 888.2900 3527.2200 891.0900 ;
      RECT 3294.6200 888.2900 3513.2600 888.3900 ;
      RECT 3285.4600 888.2900 3286.7600 891.0900 ;
      RECT 3054.1600 888.2900 3272.8000 888.3900 ;
      RECT 3045.0000 888.2900 3046.3000 891.0900 ;
      RECT 2813.7000 888.2900 3032.3400 888.3900 ;
      RECT 2804.5400 888.2900 2805.8400 891.0900 ;
      RECT 2573.2400 888.2900 2791.8800 888.3900 ;
      RECT 2564.0800 888.2900 2565.3800 891.0900 ;
      RECT 2332.7800 888.2900 2551.4200 888.3900 ;
      RECT 2323.6200 888.2900 2324.9200 891.0900 ;
      RECT 2092.3200 888.2900 2310.9600 888.3900 ;
      RECT 2083.1600 888.2900 2084.4600 891.0900 ;
      RECT 1851.8600 888.2900 2070.5000 888.3900 ;
      RECT 1842.7000 888.2900 1844.0000 891.0900 ;
      RECT 1611.4000 888.2900 1830.0400 888.3900 ;
      RECT 1602.2400 888.2900 1603.5400 891.0900 ;
      RECT 1370.9400 888.2900 1589.5800 888.3900 ;
      RECT 1361.7800 888.2900 1363.0800 891.0900 ;
      RECT 1130.4800 888.2900 1349.1200 888.3900 ;
      RECT 1121.3200 888.2900 1122.6200 891.0900 ;
      RECT 890.0200 888.2900 1108.6600 888.3900 ;
      RECT 880.8600 888.2900 882.1600 891.0900 ;
      RECT 649.5600 888.2900 868.2000 888.3900 ;
      RECT 640.4000 888.2900 641.7000 891.0900 ;
      RECT 409.1000 888.2900 627.7400 888.3900 ;
      RECT 399.9400 888.2900 401.2400 891.0900 ;
      RECT 168.6400 888.2900 387.2800 888.3900 ;
      RECT 159.3800 888.2900 160.6800 891.0900 ;
      RECT 3776.3800 884.4600 3777.7800 889.2900 ;
      RECT 3770.3800 884.4600 3773.7800 1118.9000 ;
      RECT 3816.2800 882.4600 3817.6800 891.7900 ;
      RECT 3780.3800 882.4600 3813.6800 889.2900 ;
      RECT 3756.3200 882.4600 3763.7800 895.4900 ;
      RECT 3529.9200 882.4600 3753.7200 888.2900 ;
      RECT 3515.8600 882.4600 3523.3200 895.4900 ;
      RECT 3289.4600 882.4600 3513.2600 888.2900 ;
      RECT 3275.4000 882.4600 3282.8600 895.4900 ;
      RECT 3049.0000 882.4600 3272.8000 888.2900 ;
      RECT 3034.9400 882.4600 3042.4000 895.4900 ;
      RECT 2808.5400 882.4600 3032.3400 888.2900 ;
      RECT 2794.4800 882.4600 2801.9400 895.4900 ;
      RECT 2568.0800 882.4600 2791.8800 888.2900 ;
      RECT 2554.0200 882.4600 2561.4800 895.4900 ;
      RECT 2327.6200 882.4600 2551.4200 888.2900 ;
      RECT 2313.5600 882.4600 2321.0200 895.4900 ;
      RECT 2087.1600 882.4600 2310.9600 888.2900 ;
      RECT 2073.1000 882.4600 2080.5600 895.4900 ;
      RECT 1846.7000 882.4600 2070.5000 888.2900 ;
      RECT 1832.6400 882.4600 1840.1000 895.4900 ;
      RECT 1606.2400 882.4600 1830.0400 888.2900 ;
      RECT 1592.1800 882.4600 1599.6400 895.4900 ;
      RECT 1365.7800 882.4600 1589.5800 888.2900 ;
      RECT 1351.7200 882.4600 1359.1800 895.4900 ;
      RECT 1125.3200 882.4600 1349.1200 888.2900 ;
      RECT 1111.2600 882.4600 1118.7200 895.4900 ;
      RECT 884.8600 882.4600 1108.6600 888.2900 ;
      RECT 870.8000 882.4600 878.2600 895.4900 ;
      RECT 644.4000 882.4600 868.2000 888.2900 ;
      RECT 630.3400 882.4600 637.8000 895.4900 ;
      RECT 403.9400 882.4600 627.7400 888.2900 ;
      RECT 389.8800 882.4600 397.3400 895.4900 ;
      RECT 163.3800 882.4600 387.2800 888.2900 ;
      RECT 3820.2800 878.4600 3917.8400 1118.9000 ;
      RECT 3780.3800 878.4600 3817.6800 882.4600 ;
      RECT 3770.3800 878.4600 3777.7800 884.4600 ;
      RECT 3770.3800 869.0600 3917.8400 878.4600 ;
      RECT 3529.9200 645.6500 3763.7800 882.4600 ;
      RECT 3289.4600 645.6500 3523.3200 882.4600 ;
      RECT 3049.0000 645.6500 3282.8600 882.4600 ;
      RECT 2808.5400 645.6500 3042.4000 882.4600 ;
      RECT 2568.0800 645.6500 2801.9400 882.4600 ;
      RECT 2327.6200 645.6500 2561.4800 882.4600 ;
      RECT 2087.1600 645.6500 2321.0200 882.4600 ;
      RECT 1846.7000 645.6500 2080.5600 882.4600 ;
      RECT 1606.2400 645.6500 1840.1000 882.4600 ;
      RECT 1365.7800 645.6500 1599.6400 882.4600 ;
      RECT 1125.3200 645.6500 1359.1800 882.4600 ;
      RECT 884.8600 645.6500 1118.7200 882.4600 ;
      RECT 644.4000 645.6500 878.2600 882.4600 ;
      RECT 403.9400 645.6500 637.8000 882.4600 ;
      RECT 163.3800 645.6500 397.3400 882.4600 ;
      RECT 159.3800 644.5100 160.7800 888.2900 ;
      RECT 123.4800 644.5100 156.7800 889.6500 ;
      RECT 123.4800 644.4100 150.4400 644.5100 ;
      RECT 3816.2800 644.2500 3817.6800 869.0600 ;
      RECT 3780.3800 644.2500 3813.6800 869.0600 ;
      RECT 3780.3800 644.1500 3807.3400 644.2500 ;
      RECT 123.4800 642.3100 149.7900 644.4100 ;
      RECT 159.4800 642.2100 160.7800 644.5100 ;
      RECT 123.4800 642.2100 150.4400 642.3100 ;
      RECT 3780.3800 642.0500 3806.6900 644.1500 ;
      RECT 3816.3800 641.9500 3817.6800 644.2500 ;
      RECT 3780.3800 641.9500 3807.3400 642.0500 ;
      RECT 123.4800 641.9100 156.7800 642.2100 ;
      RECT 3780.3800 641.7500 3813.6800 641.9500 ;
      RECT 3776.3800 641.7500 3777.7800 869.0600 ;
      RECT 3784.2200 641.6500 3813.6800 641.7500 ;
      RECT 3529.9200 641.2500 3753.7200 645.6500 ;
      RECT 3525.9200 641.2500 3527.3200 888.2900 ;
      RECT 3289.4600 641.2500 3513.2600 645.6500 ;
      RECT 3285.4600 641.2500 3286.8600 888.2900 ;
      RECT 3049.0000 641.2500 3272.8000 645.6500 ;
      RECT 3045.0000 641.2500 3046.4000 888.2900 ;
      RECT 2808.5400 641.2500 3032.3400 645.6500 ;
      RECT 2804.5400 641.2500 2805.9400 888.2900 ;
      RECT 2568.0800 641.2500 2791.8800 645.6500 ;
      RECT 2564.0800 641.2500 2565.4800 888.2900 ;
      RECT 2327.6200 641.2500 2551.4200 645.6500 ;
      RECT 2323.6200 641.2500 2325.0200 888.2900 ;
      RECT 2087.1600 641.2500 2310.9600 645.6500 ;
      RECT 2083.1600 641.2500 2084.5600 888.2900 ;
      RECT 1846.7000 641.2500 2070.5000 645.6500 ;
      RECT 1842.7000 641.2500 1844.1000 888.2900 ;
      RECT 1606.2400 641.2500 1830.0400 645.6500 ;
      RECT 1602.2400 641.2500 1603.6400 888.2900 ;
      RECT 1365.7800 641.2500 1589.5800 645.6500 ;
      RECT 1361.7800 641.2500 1363.1800 888.2900 ;
      RECT 1125.3200 641.2500 1349.1200 645.6500 ;
      RECT 1121.3200 641.2500 1122.7200 888.2900 ;
      RECT 884.8600 641.2500 1108.6600 645.6500 ;
      RECT 880.8600 641.2500 882.2600 888.2900 ;
      RECT 644.4000 641.2500 868.2000 645.6500 ;
      RECT 640.4000 641.2500 641.8000 888.2900 ;
      RECT 403.9400 641.2500 627.7400 645.6500 ;
      RECT 399.9400 641.2500 401.3400 888.2900 ;
      RECT 163.3800 641.2500 387.2800 645.6500 ;
      RECT 159.3800 641.2500 160.7800 642.2100 ;
      RECT 3535.0800 641.1500 3753.7200 641.2500 ;
      RECT 3294.6200 641.1500 3513.2600 641.2500 ;
      RECT 3054.1600 641.1500 3272.8000 641.2500 ;
      RECT 2813.7000 641.1500 3032.3400 641.2500 ;
      RECT 2573.2400 641.1500 2791.8800 641.2500 ;
      RECT 2332.7800 641.1500 2551.4200 641.2500 ;
      RECT 2092.3200 641.1500 2310.9600 641.2500 ;
      RECT 1851.8600 641.1500 2070.5000 641.2500 ;
      RECT 1611.4000 641.1500 1830.0400 641.2500 ;
      RECT 1370.9400 641.1500 1589.5800 641.2500 ;
      RECT 1130.4800 641.1500 1349.1200 641.2500 ;
      RECT 890.0200 641.1500 1108.6600 641.2500 ;
      RECT 649.5600 641.1500 868.2000 641.2500 ;
      RECT 409.1000 641.1500 627.7400 641.2500 ;
      RECT 168.6400 641.1500 387.2800 641.2500 ;
      RECT 156.3100 639.8100 156.7800 641.9100 ;
      RECT 123.4800 639.8100 151.7050 641.9100 ;
      RECT 3784.8700 639.5500 3813.6800 641.6500 ;
      RECT 3784.2200 639.4500 3813.6800 639.5500 ;
      RECT 3776.3800 639.4500 3777.6800 641.7500 ;
      RECT 3536.4800 638.5500 3753.7200 641.1500 ;
      RECT 3296.0200 638.5500 3513.2600 641.1500 ;
      RECT 3055.5600 638.5500 3272.8000 641.1500 ;
      RECT 2815.1000 638.5500 3032.3400 641.1500 ;
      RECT 2574.6400 638.5500 2791.8800 641.1500 ;
      RECT 2334.1800 638.5500 2551.4200 641.1500 ;
      RECT 2093.7200 638.5500 2310.9600 641.1500 ;
      RECT 1853.2600 638.5500 2070.5000 641.1500 ;
      RECT 1612.8000 638.5500 1830.0400 641.1500 ;
      RECT 1372.3400 638.5500 1589.5800 641.1500 ;
      RECT 1131.8800 638.5500 1349.1200 641.1500 ;
      RECT 891.4200 638.5500 1108.6600 641.1500 ;
      RECT 650.9600 638.5500 868.2000 641.1500 ;
      RECT 410.5000 638.5500 627.7400 641.1500 ;
      RECT 170.0400 638.5500 387.2800 641.1500 ;
      RECT 3535.0800 638.4500 3753.7200 638.5500 ;
      RECT 3525.9200 638.4500 3527.2200 641.2500 ;
      RECT 3294.6200 638.4500 3513.2600 638.5500 ;
      RECT 3285.4600 638.4500 3286.7600 641.2500 ;
      RECT 3054.1600 638.4500 3272.8000 638.5500 ;
      RECT 3045.0000 638.4500 3046.3000 641.2500 ;
      RECT 2813.7000 638.4500 3032.3400 638.5500 ;
      RECT 2804.5400 638.4500 2805.8400 641.2500 ;
      RECT 2573.2400 638.4500 2791.8800 638.5500 ;
      RECT 2564.0800 638.4500 2565.3800 641.2500 ;
      RECT 2332.7800 638.4500 2551.4200 638.5500 ;
      RECT 2323.6200 638.4500 2324.9200 641.2500 ;
      RECT 2092.3200 638.4500 2310.9600 638.5500 ;
      RECT 2083.1600 638.4500 2084.4600 641.2500 ;
      RECT 1851.8600 638.4500 2070.5000 638.5500 ;
      RECT 1842.7000 638.4500 1844.0000 641.2500 ;
      RECT 1611.4000 638.4500 1830.0400 638.5500 ;
      RECT 1602.2400 638.4500 1603.5400 641.2500 ;
      RECT 1370.9400 638.4500 1589.5800 638.5500 ;
      RECT 1361.7800 638.4500 1363.0800 641.2500 ;
      RECT 1130.4800 638.4500 1349.1200 638.5500 ;
      RECT 1121.3200 638.4500 1122.6200 641.2500 ;
      RECT 890.0200 638.4500 1108.6600 638.5500 ;
      RECT 880.8600 638.4500 882.1600 641.2500 ;
      RECT 649.5600 638.4500 868.2000 638.5500 ;
      RECT 640.4000 638.4500 641.7000 641.2500 ;
      RECT 409.1000 638.4500 627.7400 638.5500 ;
      RECT 399.9400 638.4500 401.2400 641.2500 ;
      RECT 168.6400 638.4500 387.2800 638.5500 ;
      RECT 159.3800 638.4500 160.6800 641.2500 ;
      RECT 3776.3800 634.6200 3777.7800 639.4500 ;
      RECT 3770.3800 634.6200 3773.7800 869.0600 ;
      RECT 3816.2800 632.6200 3817.6800 641.9500 ;
      RECT 3780.3800 632.6200 3813.6800 639.4500 ;
      RECT 3756.3200 632.6200 3763.7800 645.6500 ;
      RECT 3529.9200 632.6200 3753.7200 638.4500 ;
      RECT 3515.8600 632.6200 3523.3200 645.6500 ;
      RECT 3289.4600 632.6200 3513.2600 638.4500 ;
      RECT 3275.4000 632.6200 3282.8600 645.6500 ;
      RECT 3049.0000 632.6200 3272.8000 638.4500 ;
      RECT 3034.9400 632.6200 3042.4000 645.6500 ;
      RECT 2808.5400 632.6200 3032.3400 638.4500 ;
      RECT 2794.4800 632.6200 2801.9400 645.6500 ;
      RECT 2568.0800 632.6200 2791.8800 638.4500 ;
      RECT 2554.0200 632.6200 2561.4800 645.6500 ;
      RECT 2327.6200 632.6200 2551.4200 638.4500 ;
      RECT 2313.5600 632.6200 2321.0200 645.6500 ;
      RECT 2087.1600 632.6200 2310.9600 638.4500 ;
      RECT 2073.1000 632.6200 2080.5600 645.6500 ;
      RECT 1846.7000 632.6200 2070.5000 638.4500 ;
      RECT 1832.6400 632.6200 1840.1000 645.6500 ;
      RECT 1606.2400 632.6200 1830.0400 638.4500 ;
      RECT 1592.1800 632.6200 1599.6400 645.6500 ;
      RECT 1365.7800 632.6200 1589.5800 638.4500 ;
      RECT 1351.7200 632.6200 1359.1800 645.6500 ;
      RECT 1125.3200 632.6200 1349.1200 638.4500 ;
      RECT 1111.2600 632.6200 1118.7200 645.6500 ;
      RECT 884.8600 632.6200 1108.6600 638.4500 ;
      RECT 870.8000 632.6200 878.2600 645.6500 ;
      RECT 644.4000 632.6200 868.2000 638.4500 ;
      RECT 630.3400 632.6200 637.8000 645.6500 ;
      RECT 403.9400 632.6200 627.7400 638.4500 ;
      RECT 389.8800 632.6200 397.3400 645.6500 ;
      RECT 163.3800 632.6200 387.2800 638.4500 ;
      RECT 3820.2800 628.6200 3917.8400 869.0600 ;
      RECT 3780.3800 628.6200 3817.6800 632.6200 ;
      RECT 3770.3800 628.6200 3777.7800 634.6200 ;
      RECT 3770.3800 619.2200 3917.8400 628.6200 ;
      RECT 3529.9200 395.8100 3763.7800 632.6200 ;
      RECT 3289.4600 395.8100 3523.3200 632.6200 ;
      RECT 3049.0000 395.8100 3282.8600 632.6200 ;
      RECT 2808.5400 395.8100 3042.4000 632.6200 ;
      RECT 2568.0800 395.8100 2801.9400 632.6200 ;
      RECT 2327.6200 395.8100 2561.4800 632.6200 ;
      RECT 2087.1600 395.8100 2321.0200 632.6200 ;
      RECT 1846.7000 395.8100 2080.5600 632.6200 ;
      RECT 1606.2400 395.8100 1840.1000 632.6200 ;
      RECT 1365.7800 395.8100 1599.6400 632.6200 ;
      RECT 1125.3200 395.8100 1359.1800 632.6200 ;
      RECT 884.8600 395.8100 1118.7200 632.6200 ;
      RECT 644.4000 395.8100 878.2600 632.6200 ;
      RECT 403.9400 395.8100 637.8000 632.6200 ;
      RECT 163.3800 395.8100 397.3400 632.6200 ;
      RECT 159.3800 394.6700 160.7800 638.4500 ;
      RECT 123.4800 394.6700 156.7800 639.8100 ;
      RECT 123.4800 394.5700 150.4400 394.6700 ;
      RECT 3816.2800 394.4100 3817.6800 619.2200 ;
      RECT 3780.3800 394.4100 3813.6800 619.2200 ;
      RECT 3780.3800 394.3100 3807.3400 394.4100 ;
      RECT 123.4800 392.4700 149.7900 394.5700 ;
      RECT 159.4800 392.3700 160.7800 394.6700 ;
      RECT 123.4800 392.3700 150.4400 392.4700 ;
      RECT 3780.3800 392.2100 3806.6900 394.3100 ;
      RECT 3816.3800 392.1100 3817.6800 394.4100 ;
      RECT 3780.3800 392.1100 3807.3400 392.2100 ;
      RECT 123.4800 392.0700 156.7800 392.3700 ;
      RECT 3780.3800 391.9100 3813.6800 392.1100 ;
      RECT 3776.3800 391.9100 3777.7800 619.2200 ;
      RECT 3784.2200 391.8100 3813.6800 391.9100 ;
      RECT 3529.9200 391.4100 3753.7200 395.8100 ;
      RECT 3525.9200 391.4100 3527.3200 638.4500 ;
      RECT 3289.4600 391.4100 3513.2600 395.8100 ;
      RECT 3285.4600 391.4100 3286.8600 638.4500 ;
      RECT 3049.0000 391.4100 3272.8000 395.8100 ;
      RECT 3045.0000 391.4100 3046.4000 638.4500 ;
      RECT 2808.5400 391.4100 3032.3400 395.8100 ;
      RECT 2804.5400 391.4100 2805.9400 638.4500 ;
      RECT 2568.0800 391.4100 2791.8800 395.8100 ;
      RECT 2564.0800 391.4100 2565.4800 638.4500 ;
      RECT 2327.6200 391.4100 2551.4200 395.8100 ;
      RECT 2323.6200 391.4100 2325.0200 638.4500 ;
      RECT 2087.1600 391.4100 2310.9600 395.8100 ;
      RECT 2083.1600 391.4100 2084.5600 638.4500 ;
      RECT 1846.7000 391.4100 2070.5000 395.8100 ;
      RECT 1842.7000 391.4100 1844.1000 638.4500 ;
      RECT 1606.2400 391.4100 1830.0400 395.8100 ;
      RECT 1602.2400 391.4100 1603.6400 638.4500 ;
      RECT 1365.7800 391.4100 1589.5800 395.8100 ;
      RECT 1361.7800 391.4100 1363.1800 638.4500 ;
      RECT 1125.3200 391.4100 1349.1200 395.8100 ;
      RECT 1121.3200 391.4100 1122.7200 638.4500 ;
      RECT 884.8600 391.4100 1108.6600 395.8100 ;
      RECT 880.8600 391.4100 882.2600 638.4500 ;
      RECT 644.4000 391.4100 868.2000 395.8100 ;
      RECT 640.4000 391.4100 641.8000 638.4500 ;
      RECT 403.9400 391.4100 627.7400 395.8100 ;
      RECT 399.9400 391.4100 401.3400 638.4500 ;
      RECT 163.3800 391.4100 387.2800 395.8100 ;
      RECT 159.3800 391.4100 160.7800 392.3700 ;
      RECT 3535.0800 391.3100 3753.7200 391.4100 ;
      RECT 3294.6200 391.3100 3513.2600 391.4100 ;
      RECT 3054.1600 391.3100 3272.8000 391.4100 ;
      RECT 2813.7000 391.3100 3032.3400 391.4100 ;
      RECT 2573.2400 391.3100 2791.8800 391.4100 ;
      RECT 2332.7800 391.3100 2551.4200 391.4100 ;
      RECT 2092.3200 391.3100 2310.9600 391.4100 ;
      RECT 1851.8600 391.3100 2070.5000 391.4100 ;
      RECT 1611.4000 391.3100 1830.0400 391.4100 ;
      RECT 1370.9400 391.3100 1589.5800 391.4100 ;
      RECT 1130.4800 391.3100 1349.1200 391.4100 ;
      RECT 890.0200 391.3100 1108.6600 391.4100 ;
      RECT 649.5600 391.3100 868.2000 391.4100 ;
      RECT 409.1000 391.3100 627.7400 391.4100 ;
      RECT 168.6400 391.3100 387.2800 391.4100 ;
      RECT 156.3100 389.9700 156.7800 392.0700 ;
      RECT 123.4800 389.9700 151.7050 392.0700 ;
      RECT 3784.8700 389.7100 3813.6800 391.8100 ;
      RECT 3784.2200 389.6100 3813.6800 389.7100 ;
      RECT 3776.3800 389.6100 3777.6800 391.9100 ;
      RECT 3536.4800 388.7100 3753.7200 391.3100 ;
      RECT 3296.0200 388.7100 3513.2600 391.3100 ;
      RECT 3055.5600 388.7100 3272.8000 391.3100 ;
      RECT 2815.1000 388.7100 3032.3400 391.3100 ;
      RECT 2574.6400 388.7100 2791.8800 391.3100 ;
      RECT 2334.1800 388.7100 2551.4200 391.3100 ;
      RECT 2093.7200 388.7100 2310.9600 391.3100 ;
      RECT 1853.2600 388.7100 2070.5000 391.3100 ;
      RECT 1612.8000 388.7100 1830.0400 391.3100 ;
      RECT 1372.3400 388.7100 1589.5800 391.3100 ;
      RECT 1131.8800 388.7100 1349.1200 391.3100 ;
      RECT 891.4200 388.7100 1108.6600 391.3100 ;
      RECT 650.9600 388.7100 868.2000 391.3100 ;
      RECT 410.5000 388.7100 627.7400 391.3100 ;
      RECT 170.0400 388.7100 387.2800 391.3100 ;
      RECT 3535.0800 388.6100 3753.7200 388.7100 ;
      RECT 3525.9200 388.6100 3527.2200 391.4100 ;
      RECT 3294.6200 388.6100 3513.2600 388.7100 ;
      RECT 3285.4600 388.6100 3286.7600 391.4100 ;
      RECT 3054.1600 388.6100 3272.8000 388.7100 ;
      RECT 3045.0000 388.6100 3046.3000 391.4100 ;
      RECT 2813.7000 388.6100 3032.3400 388.7100 ;
      RECT 2804.5400 388.6100 2805.8400 391.4100 ;
      RECT 2573.2400 388.6100 2791.8800 388.7100 ;
      RECT 2564.0800 388.6100 2565.3800 391.4100 ;
      RECT 2332.7800 388.6100 2551.4200 388.7100 ;
      RECT 2323.6200 388.6100 2324.9200 391.4100 ;
      RECT 2092.3200 388.6100 2310.9600 388.7100 ;
      RECT 2083.1600 388.6100 2084.4600 391.4100 ;
      RECT 1851.8600 388.6100 2070.5000 388.7100 ;
      RECT 1842.7000 388.6100 1844.0000 391.4100 ;
      RECT 1611.4000 388.6100 1830.0400 388.7100 ;
      RECT 1602.2400 388.6100 1603.5400 391.4100 ;
      RECT 1370.9400 388.6100 1589.5800 388.7100 ;
      RECT 1361.7800 388.6100 1363.0800 391.4100 ;
      RECT 1130.4800 388.6100 1349.1200 388.7100 ;
      RECT 1121.3200 388.6100 1122.6200 391.4100 ;
      RECT 890.0200 388.6100 1108.6600 388.7100 ;
      RECT 880.8600 388.6100 882.1600 391.4100 ;
      RECT 649.5600 388.6100 868.2000 388.7100 ;
      RECT 640.4000 388.6100 641.7000 391.4100 ;
      RECT 409.1000 388.6100 627.7400 388.7100 ;
      RECT 399.9400 388.6100 401.2400 391.4100 ;
      RECT 168.6400 388.6100 387.2800 388.7100 ;
      RECT 159.3800 388.6100 160.6800 391.4100 ;
      RECT 3776.3800 384.7800 3777.7800 389.6100 ;
      RECT 3770.3800 384.7800 3773.7800 619.2200 ;
      RECT 3816.2800 382.7800 3817.6800 392.1100 ;
      RECT 3780.3800 382.7800 3813.6800 389.6100 ;
      RECT 3756.3200 382.7800 3763.7800 395.8100 ;
      RECT 3529.9200 382.7800 3753.7200 388.6100 ;
      RECT 3515.8600 382.7800 3523.3200 395.8100 ;
      RECT 3289.4600 382.7800 3513.2600 388.6100 ;
      RECT 3275.4000 382.7800 3282.8600 395.8100 ;
      RECT 3049.0000 382.7800 3272.8000 388.6100 ;
      RECT 3034.9400 382.7800 3042.4000 395.8100 ;
      RECT 2808.5400 382.7800 3032.3400 388.6100 ;
      RECT 2794.4800 382.7800 2801.9400 395.8100 ;
      RECT 2568.0800 382.7800 2791.8800 388.6100 ;
      RECT 2554.0200 382.7800 2561.4800 395.8100 ;
      RECT 2327.6200 382.7800 2551.4200 388.6100 ;
      RECT 2313.5600 382.7800 2321.0200 395.8100 ;
      RECT 2087.1600 382.7800 2310.9600 388.6100 ;
      RECT 2073.1000 382.7800 2080.5600 395.8100 ;
      RECT 1846.7000 382.7800 2070.5000 388.6100 ;
      RECT 1832.6400 382.7800 1840.1000 395.8100 ;
      RECT 1606.2400 382.7800 1830.0400 388.6100 ;
      RECT 1592.1800 382.7800 1599.6400 395.8100 ;
      RECT 1365.7800 382.7800 1589.5800 388.6100 ;
      RECT 1351.7200 382.7800 1359.1800 395.8100 ;
      RECT 1125.3200 382.7800 1349.1200 388.6100 ;
      RECT 1111.2600 382.7800 1118.7200 395.8100 ;
      RECT 884.8600 382.7800 1108.6600 388.6100 ;
      RECT 870.8000 382.7800 878.2600 395.8100 ;
      RECT 644.4000 382.7800 868.2000 388.6100 ;
      RECT 630.3400 382.7800 637.8000 395.8100 ;
      RECT 403.9400 382.7800 627.7400 388.6100 ;
      RECT 389.8800 382.7800 397.3400 395.8100 ;
      RECT 163.3800 382.7800 387.2800 388.6100 ;
      RECT 3820.2800 378.7800 3917.8400 619.2200 ;
      RECT 3780.3800 378.7800 3817.6800 382.7800 ;
      RECT 3770.3800 378.7800 3777.7800 384.7800 ;
      RECT 3770.3800 369.3800 3917.8400 378.7800 ;
      RECT 3529.9200 145.9700 3763.7800 382.7800 ;
      RECT 3289.4600 145.9700 3523.3200 382.7800 ;
      RECT 3049.0000 145.9700 3282.8600 382.7800 ;
      RECT 2808.5400 145.9700 3042.4000 382.7800 ;
      RECT 2568.0800 145.9700 2801.9400 382.7800 ;
      RECT 2327.6200 145.9700 2561.4800 382.7800 ;
      RECT 2087.1600 145.9700 2321.0200 382.7800 ;
      RECT 1846.7000 145.9700 2080.5600 382.7800 ;
      RECT 1606.2400 145.9700 1840.1000 382.7800 ;
      RECT 1365.7800 145.9700 1599.6400 382.7800 ;
      RECT 1125.3200 145.9700 1359.1800 382.7800 ;
      RECT 884.8600 145.9700 1118.7200 382.7800 ;
      RECT 644.4000 145.9700 878.2600 382.7800 ;
      RECT 403.9400 145.9700 637.8000 382.7800 ;
      RECT 163.3800 145.9700 397.3400 382.7800 ;
      RECT 159.3800 144.8300 160.7800 388.6100 ;
      RECT 123.4800 144.8300 156.7800 389.9700 ;
      RECT 123.4800 144.7300 150.4400 144.8300 ;
      RECT 3816.2800 144.5700 3817.6800 369.3800 ;
      RECT 3780.3800 144.5700 3813.6800 369.3800 ;
      RECT 3780.3800 144.4700 3807.3400 144.5700 ;
      RECT 123.4800 142.6300 149.7900 144.7300 ;
      RECT 159.4800 142.5300 160.7800 144.8300 ;
      RECT 123.4800 142.5300 150.4400 142.6300 ;
      RECT 3780.3800 142.3700 3806.6900 144.4700 ;
      RECT 3816.3800 142.2700 3817.6800 144.5700 ;
      RECT 3780.3800 142.2700 3807.3400 142.3700 ;
      RECT 123.4800 142.2300 156.7800 142.5300 ;
      RECT 3780.3800 142.0700 3813.6800 142.2700 ;
      RECT 3776.3800 142.0700 3777.7800 369.3800 ;
      RECT 3784.2200 141.9700 3813.6800 142.0700 ;
      RECT 3529.9200 141.5700 3537.3800 145.9700 ;
      RECT 3525.9200 141.5700 3527.3200 388.6100 ;
      RECT 3289.4600 141.5700 3513.2600 145.9700 ;
      RECT 3285.4600 141.5700 3286.8600 388.6100 ;
      RECT 3049.0000 141.5700 3272.8000 145.9700 ;
      RECT 3045.0000 141.5700 3046.4000 388.6100 ;
      RECT 2808.5400 141.5700 3032.3400 145.9700 ;
      RECT 2804.5400 141.5700 2805.9400 388.6100 ;
      RECT 2568.0800 141.5700 2791.8800 145.9700 ;
      RECT 2564.0800 141.5700 2565.4800 388.6100 ;
      RECT 2327.6200 141.5700 2551.4200 145.9700 ;
      RECT 2323.6200 141.5700 2325.0200 388.6100 ;
      RECT 2087.1600 141.5700 2310.9600 145.9700 ;
      RECT 2083.1600 141.5700 2084.5600 388.6100 ;
      RECT 1846.7000 141.5700 2070.5000 145.9700 ;
      RECT 1842.7000 141.5700 1844.1000 388.6100 ;
      RECT 1606.2400 141.5700 1830.0400 145.9700 ;
      RECT 1602.2400 141.5700 1603.6400 388.6100 ;
      RECT 1365.7800 141.5700 1589.5800 145.9700 ;
      RECT 1361.7800 141.5700 1363.1800 388.6100 ;
      RECT 1125.3200 141.5700 1349.1200 145.9700 ;
      RECT 1121.3200 141.5700 1122.7200 388.6100 ;
      RECT 884.8600 141.5700 1108.6600 145.9700 ;
      RECT 880.8600 141.5700 882.2600 388.6100 ;
      RECT 644.4000 141.5700 868.2000 145.9700 ;
      RECT 640.4000 141.5700 641.8000 388.6100 ;
      RECT 403.9400 141.5700 627.7400 145.9700 ;
      RECT 399.9400 141.5700 401.3400 388.6100 ;
      RECT 163.3800 141.5700 387.2800 145.9700 ;
      RECT 159.3800 141.5700 160.7800 142.5300 ;
      RECT 3535.0800 141.4700 3537.3800 141.5700 ;
      RECT 3294.6200 141.4700 3513.2600 141.5700 ;
      RECT 3054.1600 141.4700 3272.8000 141.5700 ;
      RECT 2813.7000 141.4700 3032.3400 141.5700 ;
      RECT 2573.2400 141.4700 2791.8800 141.5700 ;
      RECT 2332.7800 141.4700 2551.4200 141.5700 ;
      RECT 2092.3200 141.4700 2310.9600 141.5700 ;
      RECT 1851.8600 141.4700 2070.5000 141.5700 ;
      RECT 1611.4000 141.4700 1830.0400 141.5700 ;
      RECT 1370.9400 141.4700 1589.5800 141.5700 ;
      RECT 1130.4800 141.4700 1349.1200 141.5700 ;
      RECT 890.0200 141.4700 1108.6600 141.5700 ;
      RECT 649.5600 141.4700 868.2000 141.5700 ;
      RECT 409.1000 141.4700 627.7400 141.5700 ;
      RECT 168.6400 141.4700 387.2800 141.5700 ;
      RECT 156.3100 140.1300 156.7800 142.2300 ;
      RECT 123.4800 140.1300 151.7050 142.2300 ;
      RECT 3784.8700 139.8700 3813.6800 141.9700 ;
      RECT 3784.2200 139.7700 3813.6800 139.8700 ;
      RECT 3776.3800 139.7700 3777.6800 142.0700 ;
      RECT 3536.4800 138.8700 3537.3800 141.4700 ;
      RECT 3296.0200 138.8700 3513.2600 141.4700 ;
      RECT 3055.5600 138.8700 3272.8000 141.4700 ;
      RECT 2815.1000 138.8700 3032.3400 141.4700 ;
      RECT 2574.6400 138.8700 2791.8800 141.4700 ;
      RECT 2334.1800 138.8700 2551.4200 141.4700 ;
      RECT 2093.7200 138.8700 2310.9600 141.4700 ;
      RECT 1853.2600 138.8700 2070.5000 141.4700 ;
      RECT 1612.8000 138.8700 1830.0400 141.4700 ;
      RECT 1372.3400 138.8700 1589.5800 141.4700 ;
      RECT 1131.8800 138.8700 1349.1200 141.4700 ;
      RECT 891.4200 138.8700 1108.6600 141.4700 ;
      RECT 650.9600 138.8700 868.2000 141.4700 ;
      RECT 410.5000 138.8700 627.7400 141.4700 ;
      RECT 170.0400 138.8700 387.2800 141.4700 ;
      RECT 3535.0800 138.7700 3537.3800 138.8700 ;
      RECT 3525.9200 138.7700 3527.2200 141.5700 ;
      RECT 3294.6200 138.7700 3513.2600 138.8700 ;
      RECT 3285.4600 138.7700 3286.7600 141.5700 ;
      RECT 3054.1600 138.7700 3272.8000 138.8700 ;
      RECT 3045.0000 138.7700 3046.3000 141.5700 ;
      RECT 2813.7000 138.7700 3032.3400 138.8700 ;
      RECT 2804.5400 138.7700 2805.8400 141.5700 ;
      RECT 2573.2400 138.7700 2791.8800 138.8700 ;
      RECT 2564.0800 138.7700 2565.3800 141.5700 ;
      RECT 2332.7800 138.7700 2551.4200 138.8700 ;
      RECT 2323.6200 138.7700 2324.9200 141.5700 ;
      RECT 2092.3200 138.7700 2310.9600 138.8700 ;
      RECT 2083.1600 138.7700 2084.4600 141.5700 ;
      RECT 1851.8600 138.7700 2070.5000 138.8700 ;
      RECT 1842.7000 138.7700 1844.0000 141.5700 ;
      RECT 1611.4000 138.7700 1830.0400 138.8700 ;
      RECT 1602.2400 138.7700 1603.5400 141.5700 ;
      RECT 1370.9400 138.7700 1589.5800 138.8700 ;
      RECT 1361.7800 138.7700 1363.0800 141.5700 ;
      RECT 1130.4800 138.7700 1349.1200 138.8700 ;
      RECT 1121.3200 138.7700 1122.6200 141.5700 ;
      RECT 890.0200 138.7700 1108.6600 138.8700 ;
      RECT 880.8600 138.7700 882.1600 141.5700 ;
      RECT 649.5600 138.7700 868.2000 138.8700 ;
      RECT 640.4000 138.7700 641.7000 141.5700 ;
      RECT 409.1000 138.7700 627.7400 138.8700 ;
      RECT 399.9400 138.7700 401.2400 141.5700 ;
      RECT 168.6400 138.7700 387.2800 138.8700 ;
      RECT 159.3800 138.7700 160.6800 141.5700 ;
      RECT 3776.3800 134.9400 3777.7800 139.7700 ;
      RECT 3770.3800 134.9400 3773.7800 369.3800 ;
      RECT 123.4800 133.2000 156.7800 140.1300 ;
      RECT 119.4800 133.2000 120.8800 3922.3600 ;
      RECT 3816.2800 132.9400 3817.6800 142.2700 ;
      RECT 3780.3800 132.9400 3813.6800 139.7700 ;
      RECT 3539.9800 132.9400 3763.7800 145.9700 ;
      RECT 3529.9200 132.9400 3537.3800 138.7700 ;
      RECT 3515.8600 132.9400 3523.3200 145.9700 ;
      RECT 3289.4600 132.9400 3513.2600 138.7700 ;
      RECT 3275.4000 132.9400 3282.8600 145.9700 ;
      RECT 3049.0000 132.9400 3272.8000 138.7700 ;
      RECT 3034.9400 132.9400 3042.4000 145.9700 ;
      RECT 2808.5400 132.9400 3032.3400 138.7700 ;
      RECT 2794.4800 132.9400 2801.9400 145.9700 ;
      RECT 2568.0800 132.9400 2791.8800 138.7700 ;
      RECT 2554.0200 132.9400 2561.4800 145.9700 ;
      RECT 2327.6200 132.9400 2551.4200 138.7700 ;
      RECT 2313.5600 132.9400 2321.0200 145.9700 ;
      RECT 2087.1600 132.9400 2310.9600 138.7700 ;
      RECT 2073.1000 132.9400 2080.5600 145.9700 ;
      RECT 1846.7000 132.9400 2070.5000 138.7700 ;
      RECT 1832.6400 132.9400 1840.1000 145.9700 ;
      RECT 1606.2400 132.9400 1830.0400 138.7700 ;
      RECT 1592.1800 132.9400 1599.6400 145.9700 ;
      RECT 1365.7800 132.9400 1589.5800 138.7700 ;
      RECT 1351.7200 132.9400 1359.1800 145.9700 ;
      RECT 1125.3200 132.9400 1349.1200 138.7700 ;
      RECT 1111.2600 132.9400 1118.7200 145.9700 ;
      RECT 884.8600 132.9400 1108.6600 138.7700 ;
      RECT 870.8000 132.9400 878.2600 145.9700 ;
      RECT 644.4000 132.9400 868.2000 138.7700 ;
      RECT 630.3400 132.9400 637.8000 145.9700 ;
      RECT 403.9400 132.9400 627.7400 138.7700 ;
      RECT 389.8800 132.9400 397.3400 145.9700 ;
      RECT 163.3800 132.9400 387.2800 138.7700 ;
      RECT 159.3800 132.9400 160.7800 138.7700 ;
      RECT 119.4800 132.9400 156.7800 133.2000 ;
      RECT 119.4800 129.2000 160.7800 132.9400 ;
      RECT 12.4000 129.2000 116.8800 3922.3600 ;
      RECT 3820.2800 128.9400 3917.8400 369.3800 ;
      RECT 3780.3800 128.9400 3817.6800 132.9400 ;
      RECT 3770.3800 128.9400 3777.7800 134.9400 ;
      RECT 163.3800 128.9400 397.3400 132.9400 ;
      RECT 12.4000 128.9400 160.7800 129.2000 ;
      RECT 12.4000 119.5400 397.3400 128.9400 ;
      RECT 3529.9200 93.3500 3763.7800 132.9400 ;
      RECT 3289.4600 93.3500 3523.3200 132.9400 ;
      RECT 3049.0000 93.3500 3282.8600 132.9400 ;
      RECT 2808.5400 93.3500 3042.4000 132.9400 ;
      RECT 2568.0800 93.3500 2801.9400 132.9400 ;
      RECT 2327.6200 93.3500 2561.4800 132.9400 ;
      RECT 2087.1600 93.3500 2321.0200 132.9400 ;
      RECT 1846.7000 93.3500 2080.5600 132.9400 ;
      RECT 1606.2400 93.3500 1840.1000 132.9400 ;
      RECT 1365.7800 93.3500 1599.6400 132.9400 ;
      RECT 1125.3200 93.3500 1359.1800 132.9400 ;
      RECT 884.8600 93.3500 1118.7200 132.9400 ;
      RECT 644.4000 93.3500 878.2600 132.9400 ;
      RECT 403.9400 93.3500 637.8000 132.9400 ;
      RECT 163.4800 93.3500 397.3400 119.5400 ;
      RECT 3756.8200 90.7500 3763.7800 93.3500 ;
      RECT 3529.9200 90.7500 3754.2200 93.3500 ;
      RECT 3516.3600 90.7500 3523.3200 93.3500 ;
      RECT 3289.4600 90.7500 3513.7600 93.3500 ;
      RECT 3275.9000 90.7500 3282.8600 93.3500 ;
      RECT 3049.0000 90.7500 3273.3000 93.3500 ;
      RECT 3035.4400 90.7500 3042.4000 93.3500 ;
      RECT 2808.5400 90.7500 3032.8400 93.3500 ;
      RECT 2794.9800 90.7500 2801.9400 93.3500 ;
      RECT 2568.0800 90.7500 2792.3800 93.3500 ;
      RECT 2554.5200 90.7500 2561.4800 93.3500 ;
      RECT 2327.6200 90.7500 2551.9200 93.3500 ;
      RECT 2314.0600 90.7500 2321.0200 93.3500 ;
      RECT 2087.1600 90.7500 2311.4600 93.3500 ;
      RECT 2073.6000 90.7500 2080.5600 93.3500 ;
      RECT 1846.7000 90.7500 2071.0000 93.3500 ;
      RECT 1833.1400 90.7500 1840.1000 93.3500 ;
      RECT 1606.2400 90.7500 1830.5400 93.3500 ;
      RECT 1592.6800 90.7500 1599.6400 93.3500 ;
      RECT 1365.7800 90.7500 1590.0800 93.3500 ;
      RECT 1352.2200 90.7500 1359.1800 93.3500 ;
      RECT 1125.3200 90.7500 1349.6200 93.3500 ;
      RECT 1111.7600 90.7500 1118.7200 93.3500 ;
      RECT 884.8600 90.7500 1109.1600 93.3500 ;
      RECT 871.3000 90.7500 878.2600 93.3500 ;
      RECT 644.4000 90.7500 868.7000 93.3500 ;
      RECT 630.8400 90.7500 637.8000 93.3500 ;
      RECT 403.9400 90.7500 628.2400 93.3500 ;
      RECT 390.3800 90.7500 397.3400 93.3500 ;
      RECT 163.4800 90.7500 387.7800 93.3500 ;
      RECT 3529.9200 90.4500 3763.7800 90.7500 ;
      RECT 3525.9200 90.4500 3527.3200 138.7700 ;
      RECT 3289.4600 90.4500 3523.3200 90.7500 ;
      RECT 3285.4600 90.4500 3286.8600 138.7700 ;
      RECT 3049.0000 90.4500 3282.8600 90.7500 ;
      RECT 3045.0000 90.4500 3046.4000 138.7700 ;
      RECT 2808.5400 90.4500 3042.4000 90.7500 ;
      RECT 2804.5400 90.4500 2805.9400 138.7700 ;
      RECT 2568.0800 90.4500 2801.9400 90.7500 ;
      RECT 2564.0800 90.4500 2565.4800 138.7700 ;
      RECT 2327.6200 90.4500 2561.4800 90.7500 ;
      RECT 2323.6200 90.4500 2325.0200 138.7700 ;
      RECT 2087.1600 90.4500 2321.0200 90.7500 ;
      RECT 2083.1600 90.4500 2084.5600 138.7700 ;
      RECT 1846.7000 90.4500 2080.5600 90.7500 ;
      RECT 1842.7000 90.4500 1844.1000 138.7700 ;
      RECT 1606.2400 90.4500 1840.1000 90.7500 ;
      RECT 1602.2400 90.4500 1603.6400 138.7700 ;
      RECT 1365.7800 90.4500 1599.6400 90.7500 ;
      RECT 1361.7800 90.4500 1363.1800 138.7700 ;
      RECT 1125.3200 90.4500 1359.1800 90.7500 ;
      RECT 1121.3200 90.4500 1122.7200 138.7700 ;
      RECT 884.8600 90.4500 1118.7200 90.7500 ;
      RECT 880.8600 90.4500 882.2600 138.7700 ;
      RECT 644.4000 90.4500 878.2600 90.7500 ;
      RECT 640.4000 90.4500 641.8000 138.7700 ;
      RECT 403.9400 90.4500 637.8000 90.7500 ;
      RECT 399.9400 90.4500 401.3400 138.7700 ;
      RECT 163.4800 90.4500 397.3400 90.7500 ;
      RECT 159.4800 90.4500 160.8800 119.5400 ;
      RECT 3535.5800 90.3500 3763.7800 90.4500 ;
      RECT 3295.1200 90.3500 3523.3200 90.4500 ;
      RECT 3054.6600 90.3500 3282.8600 90.4500 ;
      RECT 2814.2000 90.3500 3042.4000 90.4500 ;
      RECT 2573.7400 90.3500 2801.9400 90.4500 ;
      RECT 2333.2800 90.3500 2561.4800 90.4500 ;
      RECT 2092.8200 90.3500 2321.0200 90.4500 ;
      RECT 1852.3600 90.3500 2080.5600 90.4500 ;
      RECT 1611.9000 90.3500 1840.1000 90.4500 ;
      RECT 1371.4400 90.3500 1599.6400 90.4500 ;
      RECT 1130.9800 90.3500 1359.1800 90.4500 ;
      RECT 890.5200 90.3500 1118.7200 90.4500 ;
      RECT 650.0600 90.3500 878.2600 90.4500 ;
      RECT 409.6000 90.3500 637.8000 90.4500 ;
      RECT 169.1400 90.3500 397.3400 90.4500 ;
      RECT 3536.4800 87.7500 3763.7800 90.3500 ;
      RECT 3296.0200 87.7500 3523.3200 90.3500 ;
      RECT 3055.5600 87.7500 3282.8600 90.3500 ;
      RECT 2815.1000 87.7500 3042.4000 90.3500 ;
      RECT 2574.6400 87.7500 2801.9400 90.3500 ;
      RECT 2334.1800 87.7500 2561.4800 90.3500 ;
      RECT 2093.7200 87.7500 2321.0200 90.3500 ;
      RECT 1853.2600 87.7500 2080.5600 90.3500 ;
      RECT 1612.8000 87.7500 1840.1000 90.3500 ;
      RECT 1372.3400 87.7500 1599.6400 90.3500 ;
      RECT 1131.8800 87.7500 1359.1800 90.3500 ;
      RECT 891.4200 87.7500 1118.7200 90.3500 ;
      RECT 650.9600 87.7500 878.2600 90.3500 ;
      RECT 410.5000 87.7500 637.8000 90.3500 ;
      RECT 170.0400 87.7500 397.3400 90.3500 ;
      RECT 3535.5800 87.6500 3763.7800 87.7500 ;
      RECT 3525.9200 87.6500 3527.2200 90.4500 ;
      RECT 3295.1200 87.6500 3523.3200 87.7500 ;
      RECT 3285.4600 87.6500 3286.7600 90.4500 ;
      RECT 3054.6600 87.6500 3282.8600 87.7500 ;
      RECT 3045.0000 87.6500 3046.3000 90.4500 ;
      RECT 2814.2000 87.6500 3042.4000 87.7500 ;
      RECT 2804.5400 87.6500 2805.8400 90.4500 ;
      RECT 2573.7400 87.6500 2801.9400 87.7500 ;
      RECT 2564.0800 87.6500 2565.3800 90.4500 ;
      RECT 2333.2800 87.6500 2561.4800 87.7500 ;
      RECT 2323.6200 87.6500 2324.9200 90.4500 ;
      RECT 2092.8200 87.6500 2321.0200 87.7500 ;
      RECT 2083.1600 87.6500 2084.4600 90.4500 ;
      RECT 1852.3600 87.6500 2080.5600 87.7500 ;
      RECT 1842.7000 87.6500 1844.0000 90.4500 ;
      RECT 1611.9000 87.6500 1840.1000 87.7500 ;
      RECT 1602.2400 87.6500 1603.5400 90.4500 ;
      RECT 1371.4400 87.6500 1599.6400 87.7500 ;
      RECT 1361.7800 87.6500 1363.0800 90.4500 ;
      RECT 1130.9800 87.6500 1359.1800 87.7500 ;
      RECT 1121.3200 87.6500 1122.6200 90.4500 ;
      RECT 890.5200 87.6500 1118.7200 87.7500 ;
      RECT 880.8600 87.6500 882.1600 90.4500 ;
      RECT 650.0600 87.6500 878.2600 87.7500 ;
      RECT 640.4000 87.6500 641.7000 90.4500 ;
      RECT 409.6000 87.6500 637.8000 87.7500 ;
      RECT 399.9400 87.6500 401.2400 90.4500 ;
      RECT 169.1400 87.6500 397.3400 87.7500 ;
      RECT 159.4800 87.6500 160.7800 90.4500 ;
      RECT 3766.3800 82.6800 3767.7800 3922.3600 ;
      RECT 3529.9200 82.6800 3763.7800 87.6500 ;
      RECT 3525.9200 82.6800 3527.3200 87.6500 ;
      RECT 3289.4600 82.6800 3523.3200 87.6500 ;
      RECT 3285.4600 82.6800 3286.8600 87.6500 ;
      RECT 3049.0000 82.6800 3282.8600 87.6500 ;
      RECT 3045.0000 82.6800 3046.4000 87.6500 ;
      RECT 2808.5400 82.6800 3042.4000 87.6500 ;
      RECT 2804.5400 82.6800 2805.9400 87.6500 ;
      RECT 2568.0800 82.6800 2801.9400 87.6500 ;
      RECT 2564.0800 82.6800 2565.4800 87.6500 ;
      RECT 2327.6200 82.6800 2561.4800 87.6500 ;
      RECT 2323.6200 82.6800 2325.0200 87.6500 ;
      RECT 2087.1600 82.6800 2321.0200 87.6500 ;
      RECT 2083.1600 82.6800 2084.5600 87.6500 ;
      RECT 1846.7000 82.6800 2080.5600 87.6500 ;
      RECT 1842.7000 82.6800 1844.1000 87.6500 ;
      RECT 1606.2400 82.6800 1840.1000 87.6500 ;
      RECT 1602.2400 82.6800 1603.6400 87.6500 ;
      RECT 1365.7800 82.6800 1599.6400 87.6500 ;
      RECT 1361.7800 82.6800 1363.1800 87.6500 ;
      RECT 1125.3200 82.6800 1359.1800 87.6500 ;
      RECT 1121.3200 82.6800 1122.7200 87.6500 ;
      RECT 884.8600 82.6800 1118.7200 87.6500 ;
      RECT 880.8600 82.6800 882.2600 87.6500 ;
      RECT 644.4000 82.6800 878.2600 87.6500 ;
      RECT 640.4000 82.6800 641.8000 87.6500 ;
      RECT 403.9400 82.6800 637.8000 87.6500 ;
      RECT 399.9400 82.6800 401.3400 87.6500 ;
      RECT 163.4800 82.6800 397.3400 87.6500 ;
      RECT 159.4800 82.6800 160.8800 87.6500 ;
      RECT 12.4000 82.6800 156.8800 119.5400 ;
      RECT 3770.3800 78.6800 3917.8400 128.9400 ;
      RECT 3529.9200 78.6800 3767.7800 82.6800 ;
      RECT 3289.4600 78.6800 3527.3200 82.6800 ;
      RECT 3049.0000 78.6800 3286.8600 82.6800 ;
      RECT 2808.5400 78.6800 3046.4000 82.6800 ;
      RECT 2568.0800 78.6800 2805.9400 82.6800 ;
      RECT 2327.6200 78.6800 2565.4800 82.6800 ;
      RECT 2087.1600 78.6800 2325.0200 82.6800 ;
      RECT 1846.7000 78.6800 2084.5600 82.6800 ;
      RECT 1606.2400 78.6800 1844.1000 82.6800 ;
      RECT 1365.7800 78.6800 1603.6400 82.6800 ;
      RECT 1125.3200 78.6800 1363.1800 82.6800 ;
      RECT 884.8600 78.6800 1122.7200 82.6800 ;
      RECT 644.4000 78.6800 882.2600 82.6800 ;
      RECT 403.9400 78.6800 641.8000 82.6800 ;
      RECT 163.4800 78.6800 401.3400 82.6800 ;
      RECT 12.4000 78.6800 160.8800 82.6800 ;
      RECT 3922.6400 7.6000 3923.8400 3922.4600 ;
      RECT 12.4000 7.6000 3917.8400 78.6800 ;
      RECT 6.4000 7.6000 7.6000 3922.4600 ;
      RECT 3928.6400 1.6000 3930.2400 3928.4600 ;
      RECT 6.4000 1.6000 3923.8400 7.6000 ;
      RECT 0.0000 1.6000 1.6000 3928.4600 ;
      RECT 0.0000 0.0000 3930.2400 1.6000 ;
    LAYER met5 ;
      RECT 0.0000 3929.6600 3930.2400 3930.0600 ;
      RECT 3929.8400 3922.4600 3930.2400 3929.6600 ;
      RECT 0.0000 3922.4600 0.4000 3929.6600 ;
      RECT 3923.8400 3916.4600 3930.2400 3922.4600 ;
      RECT 0.0000 3916.4600 6.4000 3922.4600 ;
      RECT 0.0000 3892.5100 3930.2400 3916.4600 ;
      RECT 3767.6800 3887.3100 3930.2400 3892.5100 ;
      RECT 3527.2200 3887.3100 3752.9200 3892.5100 ;
      RECT 3286.7600 3887.3100 3512.4600 3892.5100 ;
      RECT 3046.3000 3887.3100 3272.0000 3892.5100 ;
      RECT 2805.8400 3887.3100 3031.5400 3892.5100 ;
      RECT 2565.3800 3887.3100 2791.0800 3892.5100 ;
      RECT 2324.9200 3887.3100 2550.6200 3892.5100 ;
      RECT 2084.4600 3887.3100 2310.1600 3892.5100 ;
      RECT 1844.0000 3887.3100 2069.7000 3892.5100 ;
      RECT 1603.5400 3887.3100 1829.2400 3892.5100 ;
      RECT 1363.0800 3887.3100 1588.7800 3892.5100 ;
      RECT 1122.6200 3887.3100 1348.3200 3892.5100 ;
      RECT 882.1600 3887.3100 1107.8600 3892.5100 ;
      RECT 641.7000 3887.3100 867.4000 3892.5100 ;
      RECT 401.2400 3887.3100 626.9400 3892.5100 ;
      RECT 0.0000 3887.3100 386.4800 3892.5100 ;
      RECT 0.0000 3884.4400 3930.2400 3887.3100 ;
      RECT 3767.6800 3880.4400 3930.2400 3884.4400 ;
      RECT 0.0000 3879.2400 155.4800 3884.4400 ;
      RECT 3771.6800 3875.2400 3930.2400 3880.4400 ;
      RECT 0.0000 3875.2400 159.4800 3879.2400 ;
      RECT 0.0000 3874.7000 3930.2400 3875.2400 ;
      RECT 0.0000 3870.7000 6.4000 3874.7000 ;
      RECT 164.6800 3869.5000 3930.2400 3874.7000 ;
      RECT 160.6800 3865.5000 3930.2400 3869.5000 ;
      RECT 0.0000 3865.5000 0.4000 3870.7000 ;
      RECT 0.0000 3641.5400 3930.2400 3865.5000 ;
      RECT 0.0000 3641.3400 159.4800 3641.5400 ;
      RECT 0.0000 3636.5400 151.7400 3641.3400 ;
      RECT 164.6800 3636.3400 3930.2400 3641.5400 ;
      RECT 0.0000 3636.3400 159.4800 3636.5400 ;
      RECT 0.0000 3634.8600 3930.2400 3636.3400 ;
      RECT 160.6800 3634.6000 3930.2400 3634.8600 ;
      RECT 3817.5800 3630.6000 3930.2400 3634.6000 ;
      RECT 0.0000 3629.6600 0.4000 3634.8600 ;
      RECT 0.0000 3625.6600 6.4000 3629.6600 ;
      RECT 3821.5800 3625.4000 3930.2400 3630.6000 ;
      RECT 0.0000 3625.4000 159.4800 3625.6600 ;
      RECT 0.0000 3624.8600 3930.2400 3625.4000 ;
      RECT 164.6800 3619.6600 3930.2400 3624.8600 ;
      RECT 0.0000 3619.6600 115.5800 3624.8600 ;
      RECT 160.6800 3615.6600 3930.2400 3619.6600 ;
      RECT 0.0000 3615.6600 119.5800 3619.6600 ;
      RECT 0.0000 3391.7000 3930.2400 3615.6600 ;
      RECT 0.0000 3391.5000 159.4800 3391.7000 ;
      RECT 0.0000 3386.7000 151.7400 3391.5000 ;
      RECT 164.6800 3386.5000 3930.2400 3391.7000 ;
      RECT 0.0000 3386.5000 159.4800 3386.7000 ;
      RECT 0.0000 3385.0200 3930.2400 3386.5000 ;
      RECT 160.6800 3384.7600 3930.2400 3385.0200 ;
      RECT 3817.5800 3380.7600 3930.2400 3384.7600 ;
      RECT 0.0000 3379.8200 0.4000 3385.0200 ;
      RECT 0.0000 3375.8200 6.4000 3379.8200 ;
      RECT 3821.5800 3375.5600 3930.2400 3380.7600 ;
      RECT 0.0000 3375.5600 159.4800 3375.8200 ;
      RECT 0.0000 3375.0200 3930.2400 3375.5600 ;
      RECT 164.6800 3369.8200 3930.2400 3375.0200 ;
      RECT 0.0000 3369.8200 115.5800 3375.0200 ;
      RECT 160.6800 3365.8200 3930.2400 3369.8200 ;
      RECT 0.0000 3365.8200 119.5800 3369.8200 ;
      RECT 0.0000 3141.8600 3930.2400 3365.8200 ;
      RECT 0.0000 3141.6600 159.4800 3141.8600 ;
      RECT 0.0000 3136.8600 151.7400 3141.6600 ;
      RECT 164.6800 3136.6600 3930.2400 3141.8600 ;
      RECT 0.0000 3136.6600 159.4800 3136.8600 ;
      RECT 0.0000 3135.1800 3930.2400 3136.6600 ;
      RECT 160.6800 3134.9200 3930.2400 3135.1800 ;
      RECT 3817.5800 3130.9200 3930.2400 3134.9200 ;
      RECT 0.0000 3129.9800 0.4000 3135.1800 ;
      RECT 0.0000 3125.9800 6.4000 3129.9800 ;
      RECT 3821.5800 3125.7200 3930.2400 3130.9200 ;
      RECT 0.0000 3125.7200 159.4800 3125.9800 ;
      RECT 0.0000 3125.1800 3930.2400 3125.7200 ;
      RECT 164.6800 3119.9800 3930.2400 3125.1800 ;
      RECT 0.0000 3119.9800 115.5800 3125.1800 ;
      RECT 160.6800 3115.9800 3930.2400 3119.9800 ;
      RECT 0.0000 3115.9800 119.5800 3119.9800 ;
      RECT 0.0000 2892.0200 3930.2400 3115.9800 ;
      RECT 0.0000 2891.8200 159.4800 2892.0200 ;
      RECT 0.0000 2887.0200 151.7400 2891.8200 ;
      RECT 164.6800 2886.8200 3930.2400 2892.0200 ;
      RECT 0.0000 2886.8200 159.4800 2887.0200 ;
      RECT 0.0000 2885.3400 3930.2400 2886.8200 ;
      RECT 160.6800 2885.0800 3930.2400 2885.3400 ;
      RECT 3817.5800 2881.0800 3930.2400 2885.0800 ;
      RECT 0.0000 2880.1400 0.4000 2885.3400 ;
      RECT 0.0000 2876.1400 6.4000 2880.1400 ;
      RECT 3821.5800 2875.8800 3930.2400 2881.0800 ;
      RECT 0.0000 2875.8800 159.4800 2876.1400 ;
      RECT 0.0000 2875.3400 3930.2400 2875.8800 ;
      RECT 164.6800 2870.1400 3930.2400 2875.3400 ;
      RECT 0.0000 2870.1400 115.5800 2875.3400 ;
      RECT 160.6800 2866.1400 3930.2400 2870.1400 ;
      RECT 0.0000 2866.1400 119.5800 2870.1400 ;
      RECT 0.0000 2642.1800 3930.2400 2866.1400 ;
      RECT 0.0000 2641.9800 159.4800 2642.1800 ;
      RECT 0.0000 2637.1800 151.7400 2641.9800 ;
      RECT 164.6800 2636.9800 3930.2400 2642.1800 ;
      RECT 0.0000 2636.9800 159.4800 2637.1800 ;
      RECT 0.0000 2635.5000 3930.2400 2636.9800 ;
      RECT 160.6800 2635.2400 3930.2400 2635.5000 ;
      RECT 3817.5800 2631.2400 3930.2400 2635.2400 ;
      RECT 0.0000 2630.3000 0.4000 2635.5000 ;
      RECT 0.0000 2626.3000 6.4000 2630.3000 ;
      RECT 3821.5800 2626.0400 3930.2400 2631.2400 ;
      RECT 0.0000 2626.0400 159.4800 2626.3000 ;
      RECT 0.0000 2625.5000 3930.2400 2626.0400 ;
      RECT 164.6800 2620.3000 3930.2400 2625.5000 ;
      RECT 0.0000 2620.3000 115.5800 2625.5000 ;
      RECT 160.6800 2616.3000 3930.2400 2620.3000 ;
      RECT 0.0000 2616.3000 119.5800 2620.3000 ;
      RECT 0.0000 2392.3400 3930.2400 2616.3000 ;
      RECT 0.0000 2392.1400 159.4800 2392.3400 ;
      RECT 0.0000 2387.3400 151.7400 2392.1400 ;
      RECT 164.6800 2387.1400 3930.2400 2392.3400 ;
      RECT 0.0000 2387.1400 159.4800 2387.3400 ;
      RECT 0.0000 2385.6600 3930.2400 2387.1400 ;
      RECT 160.6800 2385.4000 3930.2400 2385.6600 ;
      RECT 3817.5800 2381.4000 3930.2400 2385.4000 ;
      RECT 0.0000 2380.4600 0.4000 2385.6600 ;
      RECT 0.0000 2376.4600 6.4000 2380.4600 ;
      RECT 3821.5800 2376.2000 3930.2400 2381.4000 ;
      RECT 0.0000 2376.2000 159.4800 2376.4600 ;
      RECT 0.0000 2375.6600 3930.2400 2376.2000 ;
      RECT 164.6800 2370.4600 3930.2400 2375.6600 ;
      RECT 0.0000 2370.4600 115.5800 2375.6600 ;
      RECT 160.6800 2366.4600 3930.2400 2370.4600 ;
      RECT 0.0000 2366.4600 119.5800 2370.4600 ;
      RECT 0.0000 2142.5000 3930.2400 2366.4600 ;
      RECT 0.0000 2142.3000 159.4800 2142.5000 ;
      RECT 0.0000 2137.5000 151.7400 2142.3000 ;
      RECT 164.6800 2137.3000 3930.2400 2142.5000 ;
      RECT 0.0000 2137.3000 159.4800 2137.5000 ;
      RECT 0.0000 2135.8200 3930.2400 2137.3000 ;
      RECT 160.6800 2135.5600 3930.2400 2135.8200 ;
      RECT 3817.5800 2131.5600 3930.2400 2135.5600 ;
      RECT 0.0000 2130.6200 0.4000 2135.8200 ;
      RECT 0.0000 2126.6200 6.4000 2130.6200 ;
      RECT 3821.5800 2126.3600 3930.2400 2131.5600 ;
      RECT 0.0000 2126.3600 159.4800 2126.6200 ;
      RECT 0.0000 2125.8200 3930.2400 2126.3600 ;
      RECT 164.6800 2120.6200 3930.2400 2125.8200 ;
      RECT 0.0000 2120.6200 115.5800 2125.8200 ;
      RECT 160.6800 2116.6200 3930.2400 2120.6200 ;
      RECT 0.0000 2116.6200 119.5800 2120.6200 ;
      RECT 0.0000 1892.6600 3930.2400 2116.6200 ;
      RECT 0.0000 1892.4600 159.4800 1892.6600 ;
      RECT 0.0000 1887.6600 151.7400 1892.4600 ;
      RECT 164.6800 1887.4600 3930.2400 1892.6600 ;
      RECT 0.0000 1887.4600 159.4800 1887.6600 ;
      RECT 0.0000 1885.9800 3930.2400 1887.4600 ;
      RECT 160.6800 1885.7200 3930.2400 1885.9800 ;
      RECT 3817.5800 1881.7200 3930.2400 1885.7200 ;
      RECT 0.0000 1880.7800 0.4000 1885.9800 ;
      RECT 0.0000 1876.7800 6.4000 1880.7800 ;
      RECT 3821.5800 1876.5200 3930.2400 1881.7200 ;
      RECT 0.0000 1876.5200 159.4800 1876.7800 ;
      RECT 0.0000 1875.9800 3930.2400 1876.5200 ;
      RECT 164.6800 1870.7800 3930.2400 1875.9800 ;
      RECT 0.0000 1870.7800 115.5800 1875.9800 ;
      RECT 160.6800 1866.7800 3930.2400 1870.7800 ;
      RECT 0.0000 1866.7800 119.5800 1870.7800 ;
      RECT 0.0000 1642.8200 3930.2400 1866.7800 ;
      RECT 0.0000 1642.6200 159.4800 1642.8200 ;
      RECT 0.0000 1637.8200 151.7400 1642.6200 ;
      RECT 164.6800 1637.6200 3930.2400 1642.8200 ;
      RECT 0.0000 1637.6200 159.4800 1637.8200 ;
      RECT 0.0000 1636.1400 3930.2400 1637.6200 ;
      RECT 160.6800 1635.8800 3930.2400 1636.1400 ;
      RECT 3817.5800 1631.8800 3930.2400 1635.8800 ;
      RECT 0.0000 1630.9400 0.4000 1636.1400 ;
      RECT 0.0000 1626.9400 6.4000 1630.9400 ;
      RECT 3821.5800 1626.6800 3930.2400 1631.8800 ;
      RECT 0.0000 1626.6800 159.4800 1626.9400 ;
      RECT 0.0000 1626.1400 3930.2400 1626.6800 ;
      RECT 164.6800 1620.9400 3930.2400 1626.1400 ;
      RECT 0.0000 1620.9400 115.5800 1626.1400 ;
      RECT 160.6800 1616.9400 3930.2400 1620.9400 ;
      RECT 0.0000 1616.9400 119.5800 1620.9400 ;
      RECT 0.0000 1392.9800 3930.2400 1616.9400 ;
      RECT 0.0000 1392.7800 159.4800 1392.9800 ;
      RECT 0.0000 1387.9800 151.7400 1392.7800 ;
      RECT 164.6800 1387.7800 3930.2400 1392.9800 ;
      RECT 0.0000 1387.7800 159.4800 1387.9800 ;
      RECT 0.0000 1386.3000 3930.2400 1387.7800 ;
      RECT 160.6800 1386.0400 3930.2400 1386.3000 ;
      RECT 3817.5800 1382.0400 3930.2400 1386.0400 ;
      RECT 0.0000 1381.1000 0.4000 1386.3000 ;
      RECT 0.0000 1377.1000 6.4000 1381.1000 ;
      RECT 3821.5800 1376.8400 3930.2400 1382.0400 ;
      RECT 0.0000 1376.8400 159.4800 1377.1000 ;
      RECT 0.0000 1376.3000 3930.2400 1376.8400 ;
      RECT 164.6800 1371.1000 3930.2400 1376.3000 ;
      RECT 0.0000 1371.1000 115.5800 1376.3000 ;
      RECT 160.6800 1367.1000 3930.2400 1371.1000 ;
      RECT 0.0000 1367.1000 119.5800 1371.1000 ;
      RECT 0.0000 1143.1400 3930.2400 1367.1000 ;
      RECT 0.0000 1142.9400 159.4800 1143.1400 ;
      RECT 0.0000 1138.1400 151.7400 1142.9400 ;
      RECT 164.6800 1137.9400 3930.2400 1143.1400 ;
      RECT 0.0000 1137.9400 159.4800 1138.1400 ;
      RECT 0.0000 1136.4600 3930.2400 1137.9400 ;
      RECT 160.6800 1136.2000 3930.2400 1136.4600 ;
      RECT 3817.5800 1132.2000 3930.2400 1136.2000 ;
      RECT 0.0000 1131.2600 0.4000 1136.4600 ;
      RECT 0.0000 1127.2600 6.4000 1131.2600 ;
      RECT 3821.5800 1127.0000 3930.2400 1132.2000 ;
      RECT 0.0000 1127.0000 159.4800 1127.2600 ;
      RECT 0.0000 1126.4600 3930.2400 1127.0000 ;
      RECT 164.6800 1121.2600 3930.2400 1126.4600 ;
      RECT 0.0000 1121.2600 115.5800 1126.4600 ;
      RECT 160.6800 1117.2600 3930.2400 1121.2600 ;
      RECT 0.0000 1117.2600 119.5800 1121.2600 ;
      RECT 0.0000 893.3000 3930.2400 1117.2600 ;
      RECT 0.0000 893.1000 159.4800 893.3000 ;
      RECT 0.0000 888.3000 151.7400 893.1000 ;
      RECT 164.6800 888.1000 3930.2400 893.3000 ;
      RECT 0.0000 888.1000 159.4800 888.3000 ;
      RECT 0.0000 886.6200 3930.2400 888.1000 ;
      RECT 160.6800 886.3600 3930.2400 886.6200 ;
      RECT 3817.5800 882.3600 3930.2400 886.3600 ;
      RECT 0.0000 881.4200 0.4000 886.6200 ;
      RECT 0.0000 877.4200 6.4000 881.4200 ;
      RECT 3821.5800 877.1600 3930.2400 882.3600 ;
      RECT 0.0000 877.1600 159.4800 877.4200 ;
      RECT 0.0000 876.6200 3930.2400 877.1600 ;
      RECT 164.6800 871.4200 3930.2400 876.6200 ;
      RECT 0.0000 871.4200 115.5800 876.6200 ;
      RECT 160.6800 867.4200 3930.2400 871.4200 ;
      RECT 0.0000 867.4200 119.5800 871.4200 ;
      RECT 0.0000 643.4600 3930.2400 867.4200 ;
      RECT 0.0000 643.2600 159.4800 643.4600 ;
      RECT 0.0000 638.4600 151.7400 643.2600 ;
      RECT 164.6800 638.2600 3930.2400 643.4600 ;
      RECT 0.0000 638.2600 159.4800 638.4600 ;
      RECT 0.0000 636.7800 3930.2400 638.2600 ;
      RECT 160.6800 636.5200 3930.2400 636.7800 ;
      RECT 3817.5800 632.5200 3930.2400 636.5200 ;
      RECT 0.0000 631.5800 0.4000 636.7800 ;
      RECT 0.0000 627.5800 6.4000 631.5800 ;
      RECT 3821.5800 627.3200 3930.2400 632.5200 ;
      RECT 0.0000 627.3200 159.4800 627.5800 ;
      RECT 0.0000 626.7800 3930.2400 627.3200 ;
      RECT 164.6800 621.5800 3930.2400 626.7800 ;
      RECT 0.0000 621.5800 115.5800 626.7800 ;
      RECT 160.6800 617.5800 3930.2400 621.5800 ;
      RECT 0.0000 617.5800 119.5800 621.5800 ;
      RECT 0.0000 393.6200 3930.2400 617.5800 ;
      RECT 0.0000 393.4200 159.4800 393.6200 ;
      RECT 0.0000 388.6200 151.7400 393.4200 ;
      RECT 164.6800 388.4200 3930.2400 393.6200 ;
      RECT 0.0000 388.4200 159.4800 388.6200 ;
      RECT 0.0000 386.9400 3930.2400 388.4200 ;
      RECT 160.6800 386.6800 3930.2400 386.9400 ;
      RECT 3817.5800 382.6800 3930.2400 386.6800 ;
      RECT 0.0000 381.7400 0.4000 386.9400 ;
      RECT 0.0000 377.7400 6.4000 381.7400 ;
      RECT 3821.5800 377.4800 3930.2400 382.6800 ;
      RECT 0.0000 377.4800 159.4800 377.7400 ;
      RECT 0.0000 376.9400 3930.2400 377.4800 ;
      RECT 164.6800 371.7400 3930.2400 376.9400 ;
      RECT 0.0000 371.7400 115.5800 376.9400 ;
      RECT 160.6800 367.7400 3930.2400 371.7400 ;
      RECT 0.0000 367.7400 119.5800 371.7400 ;
      RECT 0.0000 143.7800 3930.2400 367.7400 ;
      RECT 0.0000 143.5800 159.4800 143.7800 ;
      RECT 0.0000 138.7800 151.7400 143.5800 ;
      RECT 164.6800 138.5800 3930.2400 143.7800 ;
      RECT 0.0000 138.5800 159.4800 138.7800 ;
      RECT 0.0000 137.1000 3930.2400 138.5800 ;
      RECT 160.6800 136.8400 3930.2400 137.1000 ;
      RECT 3817.5800 132.8400 3930.2400 136.8400 ;
      RECT 0.0000 131.9000 0.4000 137.1000 ;
      RECT 0.0000 127.9000 6.4000 131.9000 ;
      RECT 3821.5800 127.6400 3930.2400 132.8400 ;
      RECT 0.0000 127.6400 159.4800 127.9000 ;
      RECT 0.0000 94.6500 3930.2400 127.6400 ;
      RECT 3767.6800 89.4500 3930.2400 94.6500 ;
      RECT 3527.2200 89.4500 3752.9200 94.6500 ;
      RECT 3286.7600 89.4500 3512.4600 94.6500 ;
      RECT 3046.3000 89.4500 3272.0000 94.6500 ;
      RECT 2805.8400 89.4500 3031.5400 94.6500 ;
      RECT 2565.3800 89.4500 2791.0800 94.6500 ;
      RECT 2324.9200 89.4500 2550.6200 94.6500 ;
      RECT 2084.4600 89.4500 2310.1600 94.6500 ;
      RECT 1844.0000 89.4500 2069.7000 94.6500 ;
      RECT 1603.5400 89.4500 1829.2400 94.6500 ;
      RECT 1363.0800 89.4500 1588.7800 94.6500 ;
      RECT 1122.6200 89.4500 1348.3200 94.6500 ;
      RECT 882.1600 89.4500 1107.8600 94.6500 ;
      RECT 641.7000 89.4500 867.4000 94.6500 ;
      RECT 401.2400 89.4500 626.9400 94.6500 ;
      RECT 0.0000 89.4500 386.4800 94.6500 ;
      RECT 0.0000 86.5800 3930.2400 89.4500 ;
      RECT 3767.6800 82.5800 3930.2400 86.5800 ;
      RECT 0.0000 81.3800 0.4000 86.5800 ;
      RECT 3771.6800 77.3800 3930.2400 82.5800 ;
      RECT 0.0000 77.3800 6.4000 81.3800 ;
      RECT 0.0000 13.6000 3930.2400 77.3800 ;
      RECT 3923.8400 7.6000 3930.2400 13.6000 ;
      RECT 0.0000 7.6000 6.4000 13.6000 ;
      RECT 3929.8400 0.4000 3930.2400 7.6000 ;
      RECT 0.0000 0.4000 0.4000 7.6000 ;
      RECT 0.0000 0.0000 3930.2400 0.4000 ;
  END
END eFPGA_top

END LIBRARY
