##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Tue Apr 20 13:36:03 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO N_term_single
  CLASS BLOCK ;
  SIZE 230.4600 BY 30.2600 ;
  FOREIGN N_term_single 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.5199 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.364 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 0.0000 19.1750 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.8628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.072 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 40.7813 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 211.259 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 0.0000 17.7950 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.6384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.118 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 22.8606 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 112.477 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 0.0000 16.4150 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.78505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.453 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 87.843 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 27.1296 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 122.377 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.33965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.929 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.4312 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.119 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 11.6514 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 57.0761 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 29.5850 0.0000 29.7550 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.0756 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.341 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 12.0563 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 55.7212 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 0.0000 28.3750 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.09105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.813 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.2824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 86.338 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 25.278 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 118.637 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 0.0000 26.9950 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.7256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.517 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 13.6283 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 65.9677 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 0.0000 26.0750 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.33965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.929 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.2054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 36.7725 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 193.697 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 0.0000 24.6950 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.49565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.289 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.9148 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.537 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 26.7593 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 123.686 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 23.1450 0.0000 23.3150 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.35705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.773 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.743 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 23.402 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 115.829 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 0.0000 21.9350 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.3968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.92 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5822 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.4337 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 20.3850 0.0000 20.5550 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.746 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.8598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 23.334 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 118.337 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 40.1650 0.0000 40.3350 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.78519 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 28.1279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 0.0000 38.9550 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.0956 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.441 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 11.0203 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 49.4559 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 37.8650 0.0000 38.0350 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.881 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.331 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 12.4129 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 60.2384 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 0.0000 36.6550 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.0558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.8169 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.503 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 35.1050 0.0000 35.2750 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.53603 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.6902 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 33.7250 0.0000 33.8950 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.7884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 68.8275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.05535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.3131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 0.0000 32.5150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.80673 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.6963 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 30.9650 0.0000 31.1350 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6724 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.325 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 1.20189 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 4.82828 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 0.0000 61.9550 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.5718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 31.3863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.494 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 0.0000 60.5750 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.87725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.385 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3808 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.867 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 2.70088 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 10.2397 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 59.0250 0.0000 59.1950 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5106 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.516 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 6.64027 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 20.6923 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 0.0000 57.8150 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.2796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.1104 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.409 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 5.22909 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 24.0714 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 0.0000 55.0550 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4056 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.954 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 5.26532 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 23.6337 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 0.0000 53.6750 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.66905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.493 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.2404 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.165 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 24.0303 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 111.853 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6484 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.205 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 6.70559 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 31.7778 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 0.0000 50.9150 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.91765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.609 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.1196 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.5205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7115 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.9697 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 49.8250 0.0000 49.9950 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.93505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.453 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.187 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 7.82707 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 36.1684 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 48.4450 0.0000 48.6150 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.68645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.337 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.7188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.304 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 42.8665 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.444 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 0.0000 47.2350 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.47265 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.909 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.5478 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 26.2418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 132.579 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 0.0000 45.8550 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.3458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 35.8496 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 187.1 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 44.3050 0.0000 44.4750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.01025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.365 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.9768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 32.7479 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.831 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 0.0000 43.0950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.96 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 21.9111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.218 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 0.0000 41.7150 0.3300 ;
    END
  END N4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.1400 0.0000 167.2800 0.4850 ;
    END
  END Ci
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.02 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 0.0000 65.6350 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.93 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 0.0000 64.2550 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.9988 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.92 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 88.0050 0.0000 88.1750 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.512 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 86.6250 0.0000 86.7950 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 0.0000 85.8750 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.1096 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.511 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 0.0000 84.4950 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 0.0000 83.1150 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 0.0000 81.7350 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER li1  ;
    ANTENNAPARTIALMETALAREA 3.52155 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER li1  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 0.0000 80.3550 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 78.8050 0.0000 78.9750 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 0.0000 77.5950 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.928 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 76.0450 0.0000 76.2150 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.24185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 74.6650 0.0000 74.8350 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.4048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.296 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 0.0000 73.9150 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.53645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.337 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3432 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.679 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.54 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.663 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.3228 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.577 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 0.0000 69.7750 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 0.0000 68.3950 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 5.2732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.292 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 109.6250 0.0000 109.7950 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.8898 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.412 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 108.2450 0.0000 108.4150 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.0924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.425 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 106.8650 0.0000 107.0350 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8692 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 105.4850 0.0000 105.6550 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.4448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.187 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 104.1050 0.0000 104.2750 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5548 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.998 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 102.7250 0.0000 102.8950 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.18365 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.569 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.5408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.63 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 101.3450 0.0000 101.5150 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7038 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.482 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9650 0.0000 100.1350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.3632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.779 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 98.5850 0.0000 98.7550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.56 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 97.6650 0.0000 97.8350 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.545 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 96.2850 0.0000 96.4550 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 94.9050 0.0000 95.0750 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1672 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.799 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 93.5250 0.0000 93.6950 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 92.1450 0.0000 92.3150 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.542 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.5955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 90.7650 0.0000 90.9350 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2484 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.205 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 89.3850 0.0000 89.5550 0.3300 ;
    END
  END S4BEG[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.0908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 26.6800 0.8000 26.9800 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 24.8500 0.8000 25.1500 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.7118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 202.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 23.0200 0.8000 23.3200 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 21.8000 0.8000 22.1000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 19.9700 0.8000 20.2700 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.928 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 18.7500 0.8000 19.0500 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.4488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 307.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 16.9200 0.8000 17.2200 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.0346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 252.272 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 15.0900 0.8000 15.3900 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.2101 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 349.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 13.8700 0.8000 14.1700 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 376.992 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 12.0400 0.8000 12.3400 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.9606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 198.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 10.8200 0.8000 11.1200 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.4817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 378.264 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 8.9900 0.8000 9.2900 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 69.6732 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 373.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 7.1600 0.8000 7.4600 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.1214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 343.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 5.9400 0.8000 6.2400 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.4534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 286.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 4.1100 0.8000 4.4100 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.2276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 215.968 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2.8900 0.8000 3.1900 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5563 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.88 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 27.6400 0.5950 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.4135 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.165 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.9400 0.5950 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6805 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 24.2400 0.5950 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.7069 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.559 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.5400 0.5950 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 164.941 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 20.8400 0.5950 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6467 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.258 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 19.1400 0.5950 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8823 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 164.398 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 17.4400 0.5950 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5563 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.88 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 15.7400 0.5950 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 14.0400 0.5950 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5249 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.4795 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.3208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.848 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 12.3400 0.5950 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6039 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.118 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 10.6400 0.5950 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5421 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 72.5655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.9338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.784 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 8.9400 0.5950 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.574 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 7.2400 0.5950 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.4611 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.404 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 5.5400 0.5950 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.7895 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.971 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 3.8400 0.5950 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.3328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.912 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 2.1400 0.5950 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.9708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 229.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 26.6800 230.4600 26.9800 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 24.8500 230.4600 25.1500 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.5918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 23.0200 230.4600 23.3200 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 21.8000 230.4600 22.1000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 19.9700 230.4600 20.2700 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.8883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 18.7500 230.4600 19.0500 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.3288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 16.9200 230.4600 17.2200 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.9146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 251.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 15.0900 230.4600 15.3900 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.1111 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.2 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 13.8700 230.4600 14.1700 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 375.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 12.0400 230.4600 12.3400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.8406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 10.8200 230.4600 11.1200 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.3617 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 377.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 8.9900 230.4600 9.2900 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 69.5532 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 372.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 7.1600 230.4600 7.4600 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 64.0014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 342.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 5.9400 230.4600 6.2400 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.3334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.856 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 4.1100 230.4600 4.4100 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.1076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 214.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 229.6600 2.8900 230.4600 3.1900 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5143 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.572 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 27.6400 230.4600 27.7800 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.3715 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 161.857 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 25.9400 230.4600 26.0800 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.7077 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 143.356 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 24.2400 230.4600 24.3800 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6663 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.258 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 22.5400 230.4600 22.6800 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9588 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 164.794 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 20.8400 230.4600 20.9800 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6369 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.11 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 19.1400 230.4600 19.2800 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8403 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 164.09 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 17.4400 230.4600 17.5800 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5143 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.572 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 15.7400 230.4600 15.8800 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6021 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.866 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 14.0400 230.4600 14.1800 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2161 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.9725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.3208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.848 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 12.3400 230.4600 12.4800 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5619 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.81 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 10.6400 230.4600 10.7800 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4465 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.9338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.784 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 8.9400 230.4600 9.0800 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.0933 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 115.322 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.574 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 7.2400 230.4600 7.3800 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.4191 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 162.096 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 5.5400 230.4600 5.6800 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.7475 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 163.663 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 3.8400 230.4600 3.9800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.3201 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 111.492 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.3328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.912 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 229.8650 2.1400 230.4600 2.2800 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.434 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 214.5200 0.0000 214.6600 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.4600 0.0000 209.6000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.434 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 204.8600 0.0000 205.0000 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7805 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 200.2600 0.0000 200.4000 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 195.6600 0.0000 195.8000 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7805 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.6000 0.0000 190.7400 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.0000 0.0000 186.1400 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 181.4000 0.0000 181.5400 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.8000 0.0000 176.9400 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.7400 0.0000 171.8800 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.366 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 162.5400 0.0000 162.6800 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.9400 0.0000 158.0800 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 152.8800 0.0000 153.0200 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 148.2800 0.0000 148.4200 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 143.6800 0.0000 143.8200 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.0800 0.0000 139.2200 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.756 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.0200 0.0000 134.1600 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.4200 0.0000 129.5600 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.8200 0.0000 124.9600 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.2200 0.0000 120.3600 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 214.0600 29.7750 214.2000 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.4600 29.7750 209.6000 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 204.4000 29.7750 204.5400 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.3400 29.7750 199.4800 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.2800 29.7750 194.4200 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 189.6800 29.7750 189.8200 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.6200 29.7750 184.7600 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.5600 29.7750 179.7000 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.5000 29.7750 174.6400 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 169.4400 29.7750 169.5800 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6193 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 164.8400 29.7750 164.9800 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.7800 29.7750 159.9200 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 154.2600 29.7750 154.4000 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 149.6600 29.7750 149.8000 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.1400 29.7750 144.2800 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4525 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.5400 29.7750 139.6800 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.4865 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.9400 29.7750 135.0800 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.4200 29.7750 129.5600 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.8200 29.7750 124.9600 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8425 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.2200 29.7750 120.3600 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
        RECT 222.9000 4.0700 224.9000 25.0000 ;
      LAYER met3 ;
        RECT 5.5600 4.0700 224.9000 6.0700 ;
        RECT 5.5600 23.0000 224.9000 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
        RECT 225.9000 1.0700 227.9000 28.0000 ;
      LAYER met3 ;
        RECT 2.5600 1.0700 227.9000 3.0700 ;
        RECT 2.5600 26.0000 227.9000 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.0000 0.5000 230.4600 30.2600 ;
      RECT 109.9650 0.0000 230.4600 0.5000 ;
      RECT 108.5850 0.0000 109.4550 0.5000 ;
      RECT 107.2050 0.0000 108.0750 0.5000 ;
      RECT 105.8250 0.0000 106.6950 0.5000 ;
      RECT 104.4450 0.0000 105.3150 0.5000 ;
      RECT 103.0650 0.0000 103.9350 0.5000 ;
      RECT 101.6850 0.0000 102.5550 0.5000 ;
      RECT 100.3050 0.0000 101.1750 0.5000 ;
      RECT 98.9250 0.0000 99.7950 0.5000 ;
      RECT 98.0050 0.0000 98.4150 0.5000 ;
      RECT 96.6250 0.0000 97.4950 0.5000 ;
      RECT 95.2450 0.0000 96.1150 0.5000 ;
      RECT 93.8650 0.0000 94.7350 0.5000 ;
      RECT 92.4850 0.0000 93.3550 0.5000 ;
      RECT 91.1050 0.0000 91.9750 0.5000 ;
      RECT 89.7250 0.0000 90.5950 0.5000 ;
      RECT 88.3450 0.0000 89.2150 0.5000 ;
      RECT 86.9650 0.0000 87.8350 0.5000 ;
      RECT 86.0450 0.0000 86.4550 0.5000 ;
      RECT 84.6650 0.0000 85.5350 0.5000 ;
      RECT 83.2850 0.0000 84.1550 0.5000 ;
      RECT 81.9050 0.0000 82.7750 0.5000 ;
      RECT 80.5250 0.0000 81.3950 0.5000 ;
      RECT 79.1450 0.0000 80.0150 0.5000 ;
      RECT 77.7650 0.0000 78.6350 0.5000 ;
      RECT 76.3850 0.0000 77.2550 0.5000 ;
      RECT 75.0050 0.0000 75.8750 0.5000 ;
      RECT 74.0850 0.0000 74.4950 0.5000 ;
      RECT 72.7050 0.0000 73.5750 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 69.9450 0.0000 70.8150 0.5000 ;
      RECT 68.5650 0.0000 69.4350 0.5000 ;
      RECT 67.1850 0.0000 68.0550 0.5000 ;
      RECT 65.8050 0.0000 66.6750 0.5000 ;
      RECT 64.4250 0.0000 65.2950 0.5000 ;
      RECT 63.0450 0.0000 63.9150 0.5000 ;
      RECT 62.1250 0.0000 62.5350 0.5000 ;
      RECT 60.7450 0.0000 61.6150 0.5000 ;
      RECT 59.3650 0.0000 60.2350 0.5000 ;
      RECT 57.9850 0.0000 58.8550 0.5000 ;
      RECT 56.6050 0.0000 57.4750 0.5000 ;
      RECT 55.2250 0.0000 56.0950 0.5000 ;
      RECT 53.8450 0.0000 54.7150 0.5000 ;
      RECT 52.4650 0.0000 53.3350 0.5000 ;
      RECT 51.0850 0.0000 51.9550 0.5000 ;
      RECT 50.1650 0.0000 50.5750 0.5000 ;
      RECT 48.7850 0.0000 49.6550 0.5000 ;
      RECT 47.4050 0.0000 48.2750 0.5000 ;
      RECT 46.0250 0.0000 46.8950 0.5000 ;
      RECT 44.6450 0.0000 45.5150 0.5000 ;
      RECT 43.2650 0.0000 44.1350 0.5000 ;
      RECT 41.8850 0.0000 42.7550 0.5000 ;
      RECT 40.5050 0.0000 41.3750 0.5000 ;
      RECT 39.1250 0.0000 39.9950 0.5000 ;
      RECT 38.2050 0.0000 38.6150 0.5000 ;
      RECT 36.8250 0.0000 37.6950 0.5000 ;
      RECT 35.4450 0.0000 36.3150 0.5000 ;
      RECT 34.0650 0.0000 34.9350 0.5000 ;
      RECT 32.6850 0.0000 33.5550 0.5000 ;
      RECT 31.3050 0.0000 32.1750 0.5000 ;
      RECT 29.9250 0.0000 30.7950 0.5000 ;
      RECT 28.5450 0.0000 29.4150 0.5000 ;
      RECT 27.1650 0.0000 28.0350 0.5000 ;
      RECT 26.2450 0.0000 26.6550 0.5000 ;
      RECT 24.8650 0.0000 25.7350 0.5000 ;
      RECT 23.4850 0.0000 24.3550 0.5000 ;
      RECT 22.1050 0.0000 22.9750 0.5000 ;
      RECT 20.7250 0.0000 21.5950 0.5000 ;
      RECT 19.3450 0.0000 20.2150 0.5000 ;
      RECT 17.9650 0.0000 18.8350 0.5000 ;
      RECT 16.5850 0.0000 17.4550 0.5000 ;
      RECT 15.6650 0.0000 16.0750 0.5000 ;
      RECT 0.0000 0.0000 15.1550 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 27.9200 230.4600 30.2600 ;
      RECT 0.7350 27.5000 229.7250 27.9200 ;
      RECT 0.0000 26.2200 230.4600 27.5000 ;
      RECT 0.7350 25.8000 229.7250 26.2200 ;
      RECT 0.0000 24.5200 230.4600 25.8000 ;
      RECT 0.7350 24.1000 229.7250 24.5200 ;
      RECT 0.0000 22.8200 230.4600 24.1000 ;
      RECT 0.7350 22.4000 229.7250 22.8200 ;
      RECT 0.0000 21.1200 230.4600 22.4000 ;
      RECT 0.7350 20.7000 229.7250 21.1200 ;
      RECT 0.0000 19.4200 230.4600 20.7000 ;
      RECT 0.7350 19.0000 229.7250 19.4200 ;
      RECT 0.0000 17.7200 230.4600 19.0000 ;
      RECT 0.7350 17.3000 229.7250 17.7200 ;
      RECT 0.0000 16.0200 230.4600 17.3000 ;
      RECT 0.7350 15.6000 229.7250 16.0200 ;
      RECT 0.0000 14.3200 230.4600 15.6000 ;
      RECT 0.7350 13.9000 229.7250 14.3200 ;
      RECT 0.0000 12.6200 230.4600 13.9000 ;
      RECT 0.7350 12.2000 229.7250 12.6200 ;
      RECT 0.0000 10.9200 230.4600 12.2000 ;
      RECT 0.7350 10.5000 229.7250 10.9200 ;
      RECT 0.0000 9.2200 230.4600 10.5000 ;
      RECT 0.7350 8.8000 229.7250 9.2200 ;
      RECT 0.0000 7.5200 230.4600 8.8000 ;
      RECT 0.7350 7.1000 229.7250 7.5200 ;
      RECT 0.0000 5.8200 230.4600 7.1000 ;
      RECT 0.7350 5.4000 229.7250 5.8200 ;
      RECT 0.0000 4.1200 230.4600 5.4000 ;
      RECT 0.7350 3.7000 229.7250 4.1200 ;
      RECT 0.0000 2.4200 230.4600 3.7000 ;
      RECT 0.7350 2.0000 229.7250 2.4200 ;
      RECT 0.0000 0.0000 230.4600 2.0000 ;
    LAYER met2 ;
      RECT 214.3400 29.6350 230.4600 30.2600 ;
      RECT 209.7400 29.6350 213.9200 30.2600 ;
      RECT 204.6800 29.6350 209.3200 30.2600 ;
      RECT 199.6200 29.6350 204.2600 30.2600 ;
      RECT 194.5600 29.6350 199.2000 30.2600 ;
      RECT 189.9600 29.6350 194.1400 30.2600 ;
      RECT 184.9000 29.6350 189.5400 30.2600 ;
      RECT 179.8400 29.6350 184.4800 30.2600 ;
      RECT 174.7800 29.6350 179.4200 30.2600 ;
      RECT 169.7200 29.6350 174.3600 30.2600 ;
      RECT 165.1200 29.6350 169.3000 30.2600 ;
      RECT 160.0600 29.6350 164.7000 30.2600 ;
      RECT 154.5400 29.6350 159.6400 30.2600 ;
      RECT 149.9400 29.6350 154.1200 30.2600 ;
      RECT 144.4200 29.6350 149.5200 30.2600 ;
      RECT 139.8200 29.6350 144.0000 30.2600 ;
      RECT 135.2200 29.6350 139.4000 30.2600 ;
      RECT 129.7000 29.6350 134.8000 30.2600 ;
      RECT 125.1000 29.6350 129.2800 30.2600 ;
      RECT 120.5000 29.6350 124.6800 30.2600 ;
      RECT 0.0000 29.6350 120.0800 30.2600 ;
      RECT 0.0000 28.1400 230.4600 29.6350 ;
      RECT 4.7000 25.1400 225.7600 28.1400 ;
      RECT 225.0400 3.9300 225.7600 25.1400 ;
      RECT 7.7000 3.9300 222.7600 25.1400 ;
      RECT 4.7000 3.9300 5.4200 25.1400 ;
      RECT 228.0400 0.9300 230.4600 28.1400 ;
      RECT 4.7000 0.9300 225.7600 3.9300 ;
      RECT 0.0000 0.9300 2.4200 28.1400 ;
      RECT 0.0000 0.6250 230.4600 0.9300 ;
      RECT 214.8000 0.0000 230.4600 0.6250 ;
      RECT 209.7400 0.0000 214.3800 0.6250 ;
      RECT 205.1400 0.0000 209.3200 0.6250 ;
      RECT 200.5400 0.0000 204.7200 0.6250 ;
      RECT 195.9400 0.0000 200.1200 0.6250 ;
      RECT 190.8800 0.0000 195.5200 0.6250 ;
      RECT 186.2800 0.0000 190.4600 0.6250 ;
      RECT 181.6800 0.0000 185.8600 0.6250 ;
      RECT 177.0800 0.0000 181.2600 0.6250 ;
      RECT 172.0200 0.0000 176.6600 0.6250 ;
      RECT 167.4200 0.0000 171.6000 0.6250 ;
      RECT 162.8200 0.0000 167.0000 0.6250 ;
      RECT 158.2200 0.0000 162.4000 0.6250 ;
      RECT 153.1600 0.0000 157.8000 0.6250 ;
      RECT 148.5600 0.0000 152.7400 0.6250 ;
      RECT 143.9600 0.0000 148.1400 0.6250 ;
      RECT 139.3600 0.0000 143.5400 0.6250 ;
      RECT 134.3000 0.0000 138.9400 0.6250 ;
      RECT 129.7000 0.0000 133.8800 0.6250 ;
      RECT 125.1000 0.0000 129.2800 0.6250 ;
      RECT 120.5000 0.0000 124.6800 0.6250 ;
      RECT 0.0000 0.0000 120.0800 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 230.4600 30.2600 ;
      RECT 228.2000 27.2800 230.4600 28.3000 ;
      RECT 0.0000 27.2800 2.2600 28.3000 ;
      RECT 228.2000 26.3800 229.3600 27.2800 ;
      RECT 1.1000 26.3800 2.2600 27.2800 ;
      RECT 228.2000 25.7000 230.4600 26.3800 ;
      RECT 0.0000 25.7000 2.2600 26.3800 ;
      RECT 0.0000 25.4500 230.4600 25.7000 ;
      RECT 1.1000 25.3000 229.3600 25.4500 ;
      RECT 225.2000 24.5500 229.3600 25.3000 ;
      RECT 1.1000 24.5500 5.2600 25.3000 ;
      RECT 225.2000 23.6200 230.4600 24.5500 ;
      RECT 0.0000 23.6200 5.2600 24.5500 ;
      RECT 225.2000 22.7200 229.3600 23.6200 ;
      RECT 1.1000 22.7200 5.2600 23.6200 ;
      RECT 225.2000 22.7000 230.4600 22.7200 ;
      RECT 0.0000 22.7000 5.2600 22.7200 ;
      RECT 0.0000 22.4000 230.4600 22.7000 ;
      RECT 1.1000 21.5000 229.3600 22.4000 ;
      RECT 0.0000 20.5700 230.4600 21.5000 ;
      RECT 1.1000 19.6700 229.3600 20.5700 ;
      RECT 0.0000 19.3500 230.4600 19.6700 ;
      RECT 1.1000 18.4500 229.3600 19.3500 ;
      RECT 0.0000 17.5200 230.4600 18.4500 ;
      RECT 1.1000 16.6200 229.3600 17.5200 ;
      RECT 0.0000 15.6900 230.4600 16.6200 ;
      RECT 1.1000 14.7900 229.3600 15.6900 ;
      RECT 0.0000 14.4700 230.4600 14.7900 ;
      RECT 1.1000 13.5700 229.3600 14.4700 ;
      RECT 0.0000 12.6400 230.4600 13.5700 ;
      RECT 1.1000 11.7400 229.3600 12.6400 ;
      RECT 0.0000 11.4200 230.4600 11.7400 ;
      RECT 1.1000 10.5200 229.3600 11.4200 ;
      RECT 0.0000 9.5900 230.4600 10.5200 ;
      RECT 1.1000 8.6900 229.3600 9.5900 ;
      RECT 0.0000 7.7600 230.4600 8.6900 ;
      RECT 1.1000 6.8600 229.3600 7.7600 ;
      RECT 0.0000 6.5400 230.4600 6.8600 ;
      RECT 1.1000 6.3700 229.3600 6.5400 ;
      RECT 225.2000 5.6400 229.3600 6.3700 ;
      RECT 1.1000 5.6400 5.2600 6.3700 ;
      RECT 225.2000 4.7100 230.4600 5.6400 ;
      RECT 0.0000 4.7100 5.2600 5.6400 ;
      RECT 225.2000 3.8100 229.3600 4.7100 ;
      RECT 1.1000 3.8100 5.2600 4.7100 ;
      RECT 225.2000 3.7700 230.4600 3.8100 ;
      RECT 0.0000 3.7700 5.2600 3.8100 ;
      RECT 0.0000 3.4900 230.4600 3.7700 ;
      RECT 1.1000 3.3700 229.3600 3.4900 ;
      RECT 228.2000 2.5900 229.3600 3.3700 ;
      RECT 1.1000 2.5900 2.2600 3.3700 ;
      RECT 228.2000 0.7700 230.4600 2.5900 ;
      RECT 0.0000 0.7700 2.2600 2.5900 ;
      RECT 0.0000 0.0000 230.4600 0.7700 ;
  END
END N_term_single

END LIBRARY
