##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Thu Apr 22 17:29:37 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LUT4AB
  CLASS BLOCK ;
  SIZE 230.4600 BY 229.8400 ;
  FOREIGN LUT4AB 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.0146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.352 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 229.5100 19.1750 229.8400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.35705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.773 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.0336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.814 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 229.5100 17.7950 229.8400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.28185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.861 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.01 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.932 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 229.5100 16.4150 229.8400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.1012 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.3545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.692 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.342 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 229.5100 15.4950 229.8400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.4398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.816 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.5850 229.5100 29.7550 229.8400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.2484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.124 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 229.5100 28.3750 229.8400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.1464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.192 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 229.5100 26.9950 229.8400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.6398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.216 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 229.5100 26.0750 229.8400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.64 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 229.5100 24.6950 229.8400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.1989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.7055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.8458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.1450 229.5100 23.3150 229.8400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9888 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.0036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.96 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 229.5100 21.9350 229.8400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 64.6914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 348.784 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.3850 229.5100 20.5550 229.8400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.825 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.3982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.873 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.1650 229.5100 40.3350 229.8400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.28225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 229.5100 38.9550 229.8400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.47 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.2355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 37.8650 229.5100 38.0350 229.8400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.606 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.9155 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.394 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 229.5100 36.6550 229.8400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 24.309 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 121.468 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.068 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.1050 229.5100 35.2750 229.8400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 25.2582 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 126.214 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.41 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.932 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.7250 229.5100 33.8950 229.8400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.0442 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.103 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 229.5100 32.5150 229.8400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 8.7532 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.729 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 30.9650 229.5100 31.1350 229.8400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.4098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 229.5100 61.9550 229.8400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.12585 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.501 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.2126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 229.5100 60.5750 229.8400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.58 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.782 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.0250 229.5100 59.1950 229.8400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.0788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 229.5100 57.8150 229.8400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 21.466 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 107.216 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 229.5100 56.4350 229.8400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.4426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 333.968 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 229.5100 55.0550 229.8400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7111 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.2348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 229.5100 53.6750 229.8400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.8188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.504 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 229.5100 52.2950 229.8400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.68385 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.981 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 22.4396 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 112.161 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 229.5100 50.9150 229.8400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.93505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.453 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.795 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 326.592 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 49.8250 229.5100 49.9950 229.8400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.58825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.045 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5545 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.9628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 48.4450 229.5100 48.6150 229.8400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.4988 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.4165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.68 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 229.5100 47.2350 229.8400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.76165 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.249 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 229.5100 45.8550 229.8400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.5756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 313.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 44.3050 229.5100 44.4750 229.8400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.0588 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.257 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 229.5100 43.0950 229.8400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.5178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 229.5100 41.7150 229.8400 ;
    END
  END N4BEG[0]
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 167.1400 229.3550 167.2800 229.8400 ;
    END
  END Co
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.95245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.297 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1152 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 47.7612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.013 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 0.0000 19.1750 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.5688 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.7295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.748 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8564 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.3684 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 0.0000 17.7950 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.35705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.773 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.6524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.1845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.3942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.574 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 21.0638 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.334545 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.8028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.752 LAYER met3  ;
    ANTENNAGATEAREA 1.485 LAYER met3  ;
    ANTENNAMAXAREACAR 31.7054 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 150.224 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.334545 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 0.0000 16.4150 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.36305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.133 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5334 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4175 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 12.9899 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 49.8131 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5595 LAYER met2  ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7912 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.4086 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.202626 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.728 LAYER met3  ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 26.3407 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.811 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.24303 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 31.0228 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 155.039 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.5578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7325 LAYER met4  ;
    ANTENNAMAXAREACAR 30.8074 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.459 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.208398 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 29.5850 0.0000 29.7550 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.64605 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.113 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.4248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 39.6749 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 193.849 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.344646 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 0.0000 28.3750 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 12.3295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.3832 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7325 LAYER met4  ;
    ANTENNAMAXAREACAR 28.9936 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.655 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.344762 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 0.0000 26.9950 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 56.4984 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 302.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 57.1502 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.438 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.50963 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 0.0000 26.0750 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.91505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.253 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.5586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7325 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5958 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 169.094 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.292698 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 0.0000 24.6950 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.0218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 35.7327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.419 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.323771 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 23.1450 0.0000 23.3150 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5661 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6115 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met1  ;
    ANTENNAMAXAREACAR 5.54397 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 20.4805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.248687 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.084 LAYER met2  ;
    ANTENNAGATEAREA 1.7325 LAYER met2  ;
    ANTENNAMAXAREACAR 6.37537 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.5694 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.248687 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 0.0000 21.9350 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.3496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 43.7966 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.954 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.560135 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 20.3850 0.0000 20.5550 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.1915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.3345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 29.3855 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.518 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.869421 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 29.921 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.999 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.922968 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 33.9947 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 142.48 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.922968 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 40.1650 0.0000 40.3350 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1344 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.2684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 LAYER met3  ;
    ANTENNAMAXAREACAR 51.9974 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.277 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.706746 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.816 LAYER met4  ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 80.2154 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.244 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.706746 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 0.0000 38.9550 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.7035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3201 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.405 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07452 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 37.8650 0.0000 38.0350 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.84285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.521 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.74 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 32.8784 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 137.847 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 0.0000 36.6550 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.93545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.0062 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4895 LAYER met4  ;
    ANTENNAMAXAREACAR 41.6897 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.215 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.818789 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 35.1050 0.0000 35.2750 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.354 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4895 LAYER met4  ;
    ANTENNAMAXAREACAR 30.5063 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 148.561 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.470633 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 33.7250 0.0000 33.8950 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6796 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.6066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4895 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2717 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.905 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.425746 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 0.0000 32.5150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.96445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.017 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.1434 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4675 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met1  ;
    ANTENNAMAXAREACAR 26.2008 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 122.442 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.318651 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5715 LAYER met2  ;
    ANTENNAGATEAREA 0.504 LAYER met2  ;
    ANTENNAMAXAREACAR 32.5335 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 153.338 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.487302 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.504 LAYER met3  ;
    ANTENNAMAXAREACAR 33.1903 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 157.767 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.0063 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.44 LAYER met4  ;
    ANTENNAGATEAREA 1.2465 LAYER met4  ;
    ANTENNAMAXAREACAR 45.229 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.102 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 30.9650 0.0000 31.1350 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.2735 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 140.725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8704 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.1312 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 104.467 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 0.0000 61.9550 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.7548 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 8.59178 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 39.6444 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 0.0000 60.5750 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.32005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.553 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.9416 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 104.671 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 30.339 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 143.484 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 59.0250 0.0000 59.1950 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.11057 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.5892 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 0.0000 57.8150 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 24.7649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 123.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 34.9328 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.525 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.83 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.113 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 28.4046 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 135.484 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 0.0000 55.0550 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.63 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.42963 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.2916 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 0.0000 53.6750 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.5485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.7812 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.5741 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.721 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 28.821 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 143.978 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 0.0000 50.9150 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3572 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.749 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 10.7838 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 35.0761 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 49.8250 0.0000 49.9950 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.10845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.657 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1269 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.5976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 276.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.5352 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 404.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 48.4450 0.0000 48.6150 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 4.46007 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 16.9522 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 0.0000 47.2350 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.87765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 30.9772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.608 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met2  ;
    ANTENNAMAXAREACAR 60.639 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 297.282 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 0.0000 45.8550 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.9265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.5314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5608 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 337.423 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.13333 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 44.3050 0.0000 44.4750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.3135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.7828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 62.4909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.052 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.598873 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 0.0000 43.0950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.1448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.6095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.3228 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.044 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met2  ;
    ANTENNAMAXAREACAR 52.0983 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 175.62 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 0.0000 41.7150 0.3300 ;
    END
  END N4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9884 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.663 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.8744 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8024 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 313.199 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.460202 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 167.6000 0.0000 167.7400 0.4850 ;
    END
  END Ci
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.3858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 67.4200 230.4600 67.5600 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 66.0600 230.4600 66.2000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 64.7000 230.4600 64.8400 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 63.0000 230.4600 63.1400 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 79.6600 230.4600 79.8000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.335 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.0606 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 77.9600 230.4600 78.1000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 76.6000 230.4600 76.7400 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.6848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 75.2400 230.4600 75.3800 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7975 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 73.5400 230.4600 73.6800 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.056 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 72.1800 230.4600 72.3200 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.2278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.352 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 70.4800 230.4600 70.6200 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.688 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 69.1200 230.4600 69.2600 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.9934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 91.5600 230.4600 91.7000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1294 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 90.2000 230.4600 90.3400 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.4838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 88.5000 230.4600 88.6400 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.687 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.989 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 87.1400 230.4600 87.2800 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 85.7800 230.4600 85.9200 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 84.0800 230.4600 84.2200 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 82.7200 230.4600 82.8600 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.1218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 81.0200 230.4600 81.1600 ;
    END
  END E2BEGb[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.609 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 109.5800 230.4600 109.7200 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1612 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 108.2200 230.4600 108.3600 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 106.8600 230.4600 107.0000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.9444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 422.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 105.1600 230.4600 105.3000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.742 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 103.8000 230.4600 103.9400 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 102.1000 230.4600 102.2400 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 100.7400 230.4600 100.8800 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.4766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 99.0400 230.4600 99.1800 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 97.6800 230.4600 97.8200 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 96.3200 230.4600 96.4600 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.689 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 491.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 94.6200 230.4600 94.7600 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 93.2600 230.4600 93.4000 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met2  ;
    ANTENNAMAXAREACAR 46.9223 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 223.062 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.805119 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.392 LAYER met3  ;
    ANTENNAGATEAREA 0.999 LAYER met3  ;
    ANTENNAMAXAREACAR 56.6681 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.507 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.845159 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3662 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.168 LAYER met4  ;
    ANTENNAGATEAREA 1.251 LAYER met4  ;
    ANTENNAMAXAREACAR 60.1583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.625 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.845159 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.4200 0.4850 67.5600 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.668 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.213 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.1404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.251 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3931 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.703 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.08042 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.0600 0.4850 66.2000 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.845 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.7822 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.756 LAYER met4  ;
    ANTENNAMAXAREACAR 67.4845 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.954762 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.7000 0.4850 64.8400 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 37.8012 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 164.319 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.8176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.768 LAYER met3  ;
    ANTENNAGATEAREA 0.504 LAYER met3  ;
    ANTENNAMAXAREACAR 82.1262 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 397.986 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.2127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 0.756 LAYER met4  ;
    ANTENNAMAXAREACAR 89.7321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2127 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 63.0000 0.4850 63.1400 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3706 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.9867 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.134949 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 79.6600 0.4850 79.8000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.9568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 32.1137 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.063 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.344646 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.9600 0.4850 78.1000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.562 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 30.5412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 159.453 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 76.6000 0.4850 76.7400 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.8426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 49.9801 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.40633 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.2400 0.4850 75.3800 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.2898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 43.5199 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.955 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.272323 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.5400 0.4850 73.6800 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.6143 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 19.6547 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.455 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 72.1800 0.4850 72.3200 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 7.63673 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.9758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.4800 0.4850 70.6200 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.5026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met4  ;
    ANTENNAMAXAREACAR 43.1387 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.352458 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 69.1200 0.4850 69.2600 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2781 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.6333 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.9798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.696 LAYER met3  ;
    ANTENNAGATEAREA 0.999 LAYER met3  ;
    ANTENNAMAXAREACAR 21.903 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.9578 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.5600 0.4850 91.7000 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.535 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 54.4144 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.935 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.568931 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.2000 0.4850 90.3400 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2332 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.786 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.5000 0.4850 88.6400 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.112 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.9438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 81.2823 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 414.154 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.666588 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.1400 0.4850 87.2800 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2465 LAYER met4  ;
    ANTENNAMAXAREACAR 70.6409 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 349.35 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.519391 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.7800 0.4850 85.9200 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.4528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7515 LAYER met3  ;
    ANTENNAMAXAREACAR 59.8168 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 277.306 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.575034 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.9788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.024 LAYER met4  ;
    ANTENNAGATEAREA 1.2465 LAYER met4  ;
    ANTENNAMAXAREACAR 73.438 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.329 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.575034 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.0800 0.4850 84.2200 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.8045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.8139 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 92.3804 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 472.465 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.7200 0.4850 82.8600 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.999 LAYER met4  ;
    ANTENNAMAXAREACAR 31.4084 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.878 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.488017 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.0200 0.4850 81.1600 ;
    END
  END E2END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.37414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.9778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.5800 0.4850 109.7200 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.557 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.2200 0.4850 108.3600 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.72579 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.5731 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.227 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.113 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.6246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7737 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 245.644 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.1600 0.4850 105.3000 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.929 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.0312 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 82.1859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 437.938 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.28539 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.2101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.1000 0.4850 102.2400 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5278 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.478 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.277 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.7566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 47.6704 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.568 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.7400 0.4850 100.8800 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.9796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 21.715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.208 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.0400 0.4850 99.1800 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.65091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.4492 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.6800 0.4850 97.8200 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.7836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 52.7821 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.362 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.3200 0.4850 96.4600 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.494 LAYER met4  ;
    ANTENNAMAXAREACAR 82.2204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.769 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.6200 0.4850 94.7600 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.6378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.494 LAYER met4  ;
    ANTENNAMAXAREACAR 115.33 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 604.3 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.1546 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.2600 0.4850 93.4000 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9412 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.6334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 367.456 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.93505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.453 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.8938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 0.0000 65.6350 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.8596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.192 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 0.0000 64.2550 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.01025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.365 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.315 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.4554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.84 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.082 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.373 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 88.0050 0.0000 88.1750 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.85725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.185 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.923 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.3916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 86.6250 0.0000 86.7950 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.10885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.3164 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.545 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 0.0000 85.8750 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.41485 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.841 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.618 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 0.0000 84.4950 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.3816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.834 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 0.0000 83.1150 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.8648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.2465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.362 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 0.0000 81.7350 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.83725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.985 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.7332 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 53.5885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 0.0000 80.3550 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.9904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 94.8745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 78.8050 0.0000 78.9750 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.95245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.297 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.016 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 0.0000 77.5950 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.3146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.952 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.0450 0.0000 76.2150 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.8306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 330.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 74.6650 0.0000 74.8350 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.41485 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.841 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.763 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 0.0000 73.9150 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.87725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.385 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.3205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.8616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.536 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.275 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.843 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 0.0000 69.7750 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 62.5788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 334.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 0.0000 68.3950 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.11225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.8158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.488 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 109.6250 0.0000 109.7950 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.9228 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.5365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.5018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.2450 0.0000 108.4150 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.28185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.861 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.9276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 106.8650 0.0000 107.0350 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.7238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.664 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.4850 0.0000 105.6550 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.8765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.7274 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.1050 0.0000 104.2750 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.7208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.7250 0.0000 102.8950 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 16.0136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.031 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 101.3450 0.0000 101.5150 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.281 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.6082 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 53.004 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9650 0.0000 100.1350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4588 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.2165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.316 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 98.5850 0.0000 98.7550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.35445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.417 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.0892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.3685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7864 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.814 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 97.6650 0.0000 97.8350 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 96.2850 0.0000 96.4550 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.8071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.2894 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 94.9050 0.0000 95.0750 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2333 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.6106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 302.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.5250 0.0000 93.6950 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.178 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 92.1450 0.0000 92.3150 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.825 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 16.2068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.997 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 90.7650 0.0000 90.9350 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.3316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 317.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 89.3850 0.0000 89.5550 0.3300 ;
    END
  END S4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.3898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 58.9488 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.801 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 229.5100 67.0150 229.8400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.2218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 66.2953 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.757603 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 229.5100 65.6350 229.8400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.51305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.133 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 58.3593 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 285.727 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.844157 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 229.5100 64.2550 229.8400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.7968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 276.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 87.6001 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 449.691 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 229.5100 62.8750 229.8400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.28225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.5486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 17.8691 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 93.0054 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 88.0050 229.5100 88.1750 229.8400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.422 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.3367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.4045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 21.879 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.222 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.2828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.312 LAYER met3  ;
    ANTENNAGATEAREA 1.2375 LAYER met3  ;
    ANTENNAMAXAREACAR 30.1883 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.919 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 86.6250 229.5100 86.7950 229.8400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.29925 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.705 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.6626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.087 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.8834 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 229.5100 85.8750 229.8400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.91505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.253 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6616 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 34.9534 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.297778 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 229.5100 84.4950 229.8400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.71025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.365 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0578 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 26.4892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 132.331 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 53.8966 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 267.825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.318 LAYER met2  ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 56.7145 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 281.82 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 229.5100 83.1150 229.8400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.825 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 22.7353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 113.491 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.7668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.598 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3562 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.4863 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 229.5100 81.7350 229.8400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.1524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.644 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 7.45826 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.2343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0415354 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 229.5100 80.3550 229.8400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.48865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.895 LAYER li1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER li1  ;
    ANTENNAMAXAREACAR 3.35172 LAYER li1  ;
    ANTENNAMAXSIDEAREACAR 3.89899 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 4.36343 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 8.8532 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.22 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.982 LAYER met2  ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 9.3897 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 78.8050 229.5100 78.9750 229.8400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.9932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.855 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 27.099 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 132.059 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0583838 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 229.5100 77.5950 229.8400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.29925 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.705 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 18.8981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.0835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 7.10081 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.2 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 76.0450 229.5100 76.2150 229.8400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.8778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 86.7952 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 445.24 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.515032 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 74.6650 229.5100 74.8350 229.8400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.58825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.045 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.2035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 21.0079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.057 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 229.5100 73.9150 229.8400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.37745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.797 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.2418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 76.6824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 229.5100 72.5350 229.8400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.8009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.2435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.1918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 34.2378 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.527 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 229.5100 71.1550 229.8400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.7326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 92.3786 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 495.102 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.94505 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 229.5100 69.7750 229.8400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.9596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 89.6965 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.898 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.680277 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 229.5100 68.3950 229.8400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.5668 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 67.7565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.188 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.86545 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.0397 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 109.6250 229.5100 109.7950 229.8400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.1464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 70.6545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.328 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.6664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.8539 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 108.2450 229.5100 108.4150 229.8400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.0688 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 95.27 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 26.3605 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 129.11 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 106.8650 229.5100 107.0350 229.8400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.6762 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 422.337 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 105.4850 229.5100 105.6550 229.8400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.4512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 141.666 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 39.2545 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 193.673 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 104.1050 229.5100 104.2750 229.8400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.93 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5643 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.306 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 102.7250 229.5100 102.8950 229.8400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.54825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.645 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.2148 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.9965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.198 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.07798 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.4 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 101.3450 229.5100 101.5150 229.8400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.4616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.271 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 15.734 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 67.1852 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 99.9650 229.5100 100.1350 229.8400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.4828 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.87421 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.7879 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 98.5850 229.5100 98.7550 229.8400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.97585 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.501 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.2524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 83.0908 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 439.03 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 97.6650 229.5100 97.8350 229.8400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.20405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.593 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.9264 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.0853 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 111.164 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 96.2850 229.5100 96.4550 229.8400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.29665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.349 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.701 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 53.4275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.47758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.5152 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 94.9050 229.5100 95.0750 229.8400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 28.8752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.668 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 61.5014 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 304.494 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 93.5250 229.5100 93.6950 229.8400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.49045 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.577 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.2956 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.3265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.8003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.5945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.1834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 96.0741 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 480.857 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 92.1450 229.5100 92.3150 229.8400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.83685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.161 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.1965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.2656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 21.2451 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.012 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 90.7650 229.5100 90.9350 229.8400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.3011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.3226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 71.6002 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 370.497 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 89.3850 229.5100 89.5550 229.8400 ;
    END
  END S4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.471 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.4800 0.4850 19.6200 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.447 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.7800 0.4850 17.9200 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.372 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.6488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.4200 0.4850 16.5600 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.9264 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.0600 0.4850 15.2000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.82 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.3800 0.4850 31.5200 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.4778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.0200 0.4850 30.1600 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.9398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.3200 0.4850 28.4600 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.1768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 26.9600 0.4850 27.1000 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.6000 0.4850 25.7400 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6851 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.461 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.9000 0.4850 24.0400 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.5884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.9200 0.4850 42.0600 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.3334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.4964 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 249.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.8600 0.4850 39.0000 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.6826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.5000 0.4850 37.6400 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.879 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.3972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.1400 0.4850 36.2800 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.6838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.4400 0.4850 34.5800 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.6736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.0800 0.4850 33.2200 ;
    END
  END W2BEGb[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.6400 0.4850 61.7800 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.807 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.5800 0.4850 58.7200 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 57.2200 0.4850 57.3600 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.5200 0.4850 55.6600 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 54.1600 0.4850 54.3000 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6258 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.66 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.4600 0.4850 52.6000 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.1000 0.4850 51.2400 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.827 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.203 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4466 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.4000 0.4850 49.5400 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.0400 0.4850 48.1800 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.362 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.7886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.9800 0.4850 45.1200 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.602 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.9776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 78.0267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.382 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.366581 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 19.4800 230.4600 19.6200 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.5728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.453 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.636111 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 17.7800 230.4600 17.9200 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.799 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.1514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.242 LAYER met4  ;
    ANTENNAMAXAREACAR 54.3692 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.880285 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 16.4200 230.4600 16.5600 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.0655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.116 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3751 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.399 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.615054 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.2128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.272 LAYER met3  ;
    ANTENNAGATEAREA 1.242 LAYER met3  ;
    ANTENNAMAXAREACAR 32.9876 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 165.045 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 15.0600 230.4600 15.2000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.44 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.4236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 38.4263 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.658 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.160673 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 31.3800 230.4600 31.5200 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.9742 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 83.322 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 443.335 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.472525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 30.0200 230.4600 30.1600 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 56.2998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 70.146 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 365.233 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 28.3200 230.4600 28.4600 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.5716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 48.7916 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 253.062 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 26.9600 230.4600 27.1000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.4198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 85.5337 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 444.07 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.239596 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 25.6000 230.4600 25.7400 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.466 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.1538 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.0121 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.704 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.0175 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.072 LAYER met4  ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 13.3038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 69.5807 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 23.9000 230.4600 24.0400 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.661 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 31.035 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.734 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.141212 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 22.5400 230.4600 22.6800 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.2568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met4  ;
    ANTENNAMAXAREACAR 54.8859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 285.776 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.168485 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 20.8400 230.4600 20.9800 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.6164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 63.0259 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 328.897 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 43.6200 230.4600 43.7600 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.6916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 56.4576 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.386 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 41.9200 230.4600 42.0600 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 40.497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 40.5600 230.4600 40.7000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3246 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 20.6055 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.408 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 38.8600 230.4600 39.0000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.736 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 55.3535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 238.377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 37.5000 230.4600 37.6400 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.2348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 28.8315 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 150.899 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 36.1400 230.4600 36.2800 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8272 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.857 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.749 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2612 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 259.891 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 34.4400 230.4600 34.5800 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.2742 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 73.3053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.337 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 33.0800 230.4600 33.2200 ;
    END
  END W2END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.449 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3577 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.8673 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 61.6400 230.4600 61.7800 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2974 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5266 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.989 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 59.9400 230.4600 60.0800 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 18.2962 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.6673 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 58.5800 230.4600 58.7200 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.765 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.4006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.2252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.169 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 57.2200 230.4600 57.3600 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.72 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.6 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 55.5200 230.4600 55.6600 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.522 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9531 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.4976 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 54.1600 230.4600 54.3000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.24593 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.3367 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 52.4600 230.4600 52.6000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 42.0897 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 202.562 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 51.1000 230.4600 51.2400 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3193 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4885 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.35529 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.3118 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 49.4000 230.4600 49.5400 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.529 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.1838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 81.5147 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 431.917 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 48.0400 230.4600 48.1800 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.577 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.01 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0541 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.505 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 46.6800 230.4600 46.8200 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.772 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1172 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.5202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 44.9800 230.4600 45.1200 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6284 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 12.0946 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 63.6197 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 114.3900 0.0000 114.6900 0.8000 ;
    END
  END UserCLK
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.9344 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.261912 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 1.0605 LAYER met3  ;
    ANTENNAMAXAREACAR 11.6862 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.0391 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.29963 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 81.5838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 437.936 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 64.7124 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 320.816 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.65283 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 214.3000 0.4850 214.4400 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.4424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 33.1023 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 147.959 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.710759 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.0723 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 369.792 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 52.7239 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 254.396 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 211.5800 0.4850 211.7200 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 122.779 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 658.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 82.0791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 395.303 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.12348 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 208.5200 0.4850 208.6600 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.702 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.941 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 62.3106 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 292.021 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.97673 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 205.4600 0.4850 205.6000 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met2  ;
    ANTENNAMAXAREACAR 27.5994 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.696 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.608586 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 27.7556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 107.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.641387 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 79.4622 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 427.552 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 66.0317 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 330.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.4000 0.4850 202.5400 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.6698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 325.717 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6045 LAYER met2  ;
    ANTENNAMAXAREACAR 49.9641 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 235.974 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.810245 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.288 LAYER met3  ;
    ANTENNAGATEAREA 3.6045 LAYER met3  ;
    ANTENNAMAXAREACAR 51.6992 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.487 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.832439 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.2326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.848 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 56.8573 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 273.236 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.832439 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 199.3400 0.4850 199.4800 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.0203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.3605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 50.4175 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 243.542 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.709434 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.3166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.296 LAYER met3  ;
    ANTENNAGATEAREA 3.9225 LAYER met3  ;
    ANTENNAMAXAREACAR 57.1266 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.564 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.709434 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 196.2800 0.4850 196.4200 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.459 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 110.556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 592.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 62.9176 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.07 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.2200 0.4850 193.3600 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.818 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3974 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.0991 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.477883 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.7256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.144 LAYER met3  ;
    ANTENNAGATEAREA 3.9225 LAYER met3  ;
    ANTENNAMAXAREACAR 41.355 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.291 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.662595 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.1600 0.4850 190.3000 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.746 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.431 LAYER met2  ;
    ANTENNAMAXAREACAR 20.5504 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.7841 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.492732 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.9348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAGATEAREA 3.6045 LAYER met3  ;
    ANTENNAMAXAREACAR 51.4394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 252.244 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.694445 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.264 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 53.8674 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.313 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 187.1000 0.4850 187.2400 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.386 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.5385 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 38.8839 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 184.0400 0.4850 184.1800 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.353 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.1579 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.327 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.248 LAYER met3  ;
    ANTENNAGATEAREA 2.9685 LAYER met3  ;
    ANTENNAMAXAREACAR 61.8428 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 297.585 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.981399 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9175 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.496 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 69.47 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.502 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 180.9800 0.4850 181.1200 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.4198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 175.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met2  ;
    ANTENNAMAXAREACAR 47.9892 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.627 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.520123 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAGATEAREA 2.6505 LAYER met3  ;
    ANTENNAMAXAREACAR 48.0881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.33 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.535214 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.008 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 50.5038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.334 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.535214 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.9200 0.4850 178.0600 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 57.3039 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 72.5537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.224 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.8600 0.4850 175.0000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met2  ;
    ANTENNAMAXAREACAR 23.3424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.6855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.505593 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.7378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.072 LAYER met3  ;
    ANTENNAGATEAREA 3.9225 LAYER met3  ;
    ANTENNAMAXAREACAR 43.5521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 209.683 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590024 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 171.8000 0.4850 171.9400 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.9725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met2  ;
    ANTENNAMAXAREACAR 24.223 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.344 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.490796 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.8729 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.784 LAYER met3  ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 29.005 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.097 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512354 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.8142 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.224 LAYER met4  ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 50.3895 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.929 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 168.7400 0.4850 168.8800 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.5505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met2  ;
    ANTENNAMAXAREACAR 40.0522 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 195.244 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.668098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.059 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.448 LAYER met3  ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 44.3955 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.659 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.689656 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2512 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.689656 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.6800 0.4850 165.8200 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met2  ;
    ANTENNAMAXAREACAR 27.1298 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.686 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.604803 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.7735 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.728 LAYER met3  ;
    ANTENNAGATEAREA 2.4915 LAYER met3  ;
    ANTENNAMAXAREACAR 72.323 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 347.453 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.898113 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 162.6200 0.4850 162.7600 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.2176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 86.5901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 421.853 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.696893 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 159.5600 0.4850 159.7000 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.7296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 45.1857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.43 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.610782 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.5000 0.4850 156.6400 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.2318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.598 LAYER met3  ;
    ANTENNAMAXAREACAR 29.8331 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 146.074 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.510969 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.1118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4 LAYER met4  ;
    ANTENNAGATEAREA 3.234 LAYER met4  ;
    ANTENNAMAXAREACAR 35.4849 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.560063 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 153.4400 0.4850 153.5800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.7283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 127.04 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.234 LAYER met2  ;
    ANTENNAMAXAREACAR 39.2049 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 171.789 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.646541 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 150.3800 0.4850 150.5200 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met2  ;
    ANTENNAMAXAREACAR 9.34507 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.0409 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.276048 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 10.3245 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.7824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.320419 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.1647 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.344 LAYER met4  ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 50.0564 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.3200 0.4850 147.4600 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 76.1418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 408.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7635 LAYER met4  ;
    ANTENNAMAXAREACAR 62.989 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 144.2600 0.4850 144.4000 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.7428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 28.9603 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.742 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.542829 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.1934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.128 LAYER met4  ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6941 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 237.246 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 141.2000 0.4850 141.3400 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.6048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 37.3639 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.542829 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAGATEAREA 2.4915 LAYER met4  ;
    ANTENNAMAXAREACAR 58.2319 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.509 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.1400 0.4850 138.2800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.993 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 219.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.1696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 33.5999 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.95 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.0800 0.4850 135.2200 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6045 LAYER met4  ;
    ANTENNAMAXAREACAR 54.8946 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.142 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.0438 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.5 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.4494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.234 LAYER met4  ;
    ANTENNAMAXAREACAR 31.8583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.082 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.630656 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.9600 0.4850 129.1000 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.234 LAYER met4  ;
    ANTENNAMAXAREACAR 26.6759 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.153 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.671278 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.9000 0.4850 126.0400 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.066 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4455 LAYER met4  ;
    ANTENNAMAXAREACAR 33.3518 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.668 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674634 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 122.8400 0.4850 122.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.5276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6045 LAYER met3  ;
    ANTENNAMAXAREACAR 42.0619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.452 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.516129 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 214.3000 230.4600 214.4400 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2793 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.08 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 211.5800 230.4600 211.7200 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 208.5200 230.4600 208.6600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.729 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 205.4600 230.4600 205.6000 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.211 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 257.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 202.4000 230.4600 202.5400 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 199.3400 230.4600 199.4800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.9788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 196.2800 230.4600 196.4200 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0872 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 193.2200 230.4600 193.3600 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.702 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.9742 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 190.1600 230.4600 190.3000 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 187.1000 230.4600 187.2400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 184.0400 230.4600 184.1800 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 180.9800 230.4600 181.1200 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 177.9200 230.4600 178.0600 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.2608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 174.8600 230.4600 175.0000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 171.8000 230.4600 171.9400 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 168.7400 230.4600 168.8800 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 165.6800 230.4600 165.8200 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.5376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 162.6200 230.4600 162.7600 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.337 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 159.5600 230.4600 159.7000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 156.5000 230.4600 156.6400 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.8628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.072 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 153.4400 230.4600 153.5800 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.1618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 150.3800 230.4600 150.5200 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.344 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 147.3200 230.4600 147.4600 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2774 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.224 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 144.2600 230.4600 144.4000 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4221 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1612 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 141.2000 230.4600 141.3400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 41.7018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 222.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 138.1400 230.4600 138.2800 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 135.0800 230.4600 135.2200 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 132.0200 230.4600 132.1600 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.577 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8684 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 128.9600 230.4600 129.1000 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 125.9000 230.4600 126.0400 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.183 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.1982 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 56.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 122.8400 230.4600 122.9800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 229.9750 120.1200 230.4600 120.2600 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.0048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 26.4803 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.402 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.660262 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 214.0600 0.0000 214.2000 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7446 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.562 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.25 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.9438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 39.3058 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.528 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695462 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.4600 0.0000 209.6000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0802 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.004 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met2  ;
    ANTENNAMAXAREACAR 25.7532 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.052 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.587477 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.128 LAYER met3  ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 28.7931 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.4968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.607333 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 29.3989 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 81.8886 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.637002 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 204.8600 0.0000 205.0000 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.883 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.2264 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 40.8015 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.043 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.807402 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 200.2600 0.0000 200.4000 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.258 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.2056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 35.2876 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.316 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.677987 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 195.6600 0.0000 195.8000 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.172 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.0594 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 31.583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.552 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.809015 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 191.0600 0.0000 191.2000 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.134 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.9186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 30.1297 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 90.8649 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.540131 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 186.0000 0.0000 186.1400 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.617 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1632 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2865 LAYER met4  ;
    ANTENNAMAXAREACAR 34.0332 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 150.171 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.994153 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 181.4000 0.0000 181.5400 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.5929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met2  ;
    ANTENNAMAXAREACAR 38.91 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 189.129 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.78805 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 176.8000 0.0000 176.9400 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.4726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.268 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.544 LAYER met2  ;
    ANTENNAMAXAREACAR 44.1204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 187.036 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.803774 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAGATEAREA 2.544 LAYER met3  ;
    ANTENNAMAXAREACAR 45.0099 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.964 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.819497 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.4718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2623 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 193.391 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.819497 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 172.2000 0.0000 172.3400 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.658 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.18 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7218 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.9491 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.659119 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 3.18 LAYER met3  ;
    ANTENNAMAXAREACAR 18.8259 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.6509 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.671698 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.4111 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.671698 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 162.5400 0.0000 162.6800 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.8305 LAYER met4  ;
    ANTENNAMAXAREACAR 26.377 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 97.1242 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.707489 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.9400 0.0000 158.0800 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.426 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.9136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 256.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2405 LAYER met4  ;
    ANTENNAMAXAREACAR 27.7638 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 108.999 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 153.3400 0.0000 153.4800 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 70.1931 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 376.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2405 LAYER met4  ;
    ANTENNAMAXAREACAR 42.2132 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 163.234 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.524686 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 148.7400 0.0000 148.8800 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.776 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.6718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2405 LAYER met4  ;
    ANTENNAMAXAREACAR 23.3935 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 88.1725 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.665407 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 144.1400 0.0000 144.2800 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.6176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2405 LAYER met4  ;
    ANTENNAMAXAREACAR 63.7374 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.77 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.794969 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 139.0800 0.0000 139.2200 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.141 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.4318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2405 LAYER met4  ;
    ANTENNAMAXAREACAR 28.7328 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 74.5702 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38863 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 134.4800 0.0000 134.6200 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.811 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.6228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2405 LAYER met4  ;
    ANTENNAMAXAREACAR 32.2473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 122.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.417765 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 129.4200 0.0000 129.5600 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.363 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 249.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.6045 LAYER met4  ;
    ANTENNAMAXAREACAR 29.8562 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.291 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.480056 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 125.2800 0.0000 125.4200 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.742 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.0996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.9225 LAYER met4  ;
    ANTENNAMAXAREACAR 16.1988 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 75.8101 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.431087 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 120.6800 0.0000 120.8200 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.6827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.3055 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 214.5200 229.3550 214.6600 229.8400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7055 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.0000 229.3550 209.1400 229.8400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.418 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 204.8600 229.3550 205.0000 229.8400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 200.2600 229.3550 200.4000 229.8400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 195.6600 229.3550 195.8000 229.8400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.8695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.6000 229.3550 190.7400 229.8400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.477 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 186.0000 229.3550 186.1400 229.8400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.483 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.13315 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.0902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.4000 229.3550 181.5400 229.8400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.784 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.6566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 176.8000 229.3550 176.9400 229.8400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.418 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.1946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 171.7400 229.3550 171.8800 229.8400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.797 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3484 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.5400 229.3550 162.6800 229.8400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.073 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.6286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 157.9400 229.3550 158.0800 229.8400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 152.8800 229.3550 153.0200 229.8400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 148.2800 229.3550 148.4200 229.8400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0565 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 143.6800 229.3550 143.8200 229.8400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.0800 229.3550 139.2200 229.8400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.0200 229.3550 134.1600 229.8400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6285 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 129.4200 229.3550 129.5600 229.8400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4705 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.8200 229.3550 124.9600 229.8400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.681 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.0406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 120.2200 229.3550 120.3600 229.8400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 190.1200 5.4300 191.7200 224.0700 ;
        RECT 160.1200 5.4300 161.7200 224.0700 ;
        RECT 130.1200 5.4300 131.7200 224.0700 ;
        RECT 100.1200 5.4300 101.7200 224.0700 ;
        RECT 70.1200 5.4300 71.7200 224.0700 ;
        RECT 40.1200 5.4300 41.7200 224.0700 ;
        RECT 221.9000 5.4300 224.9000 224.0700 ;
        RECT 5.5600 5.4300 8.5600 224.0700 ;
      LAYER met3 ;
        RECT 5.5600 5.4300 224.9000 8.4300 ;
        RECT 5.5600 221.0700 224.9000 224.0700 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 193.3200 1.4300 194.9200 228.0700 ;
        RECT 163.3200 1.4300 164.9200 228.0700 ;
        RECT 133.3200 1.4300 134.9200 228.0700 ;
        RECT 103.3200 1.4300 104.9200 228.0700 ;
        RECT 73.3200 1.4300 74.9200 228.0700 ;
        RECT 43.3200 1.4300 44.9200 228.0700 ;
        RECT 13.3200 1.4300 14.9200 228.0700 ;
        RECT 225.9000 1.4300 228.9000 228.0700 ;
        RECT 1.5600 1.4300 4.5600 228.0700 ;
      LAYER met3 ;
        RECT 1.5600 1.4300 228.9000 4.4300 ;
        RECT 1.5600 225.0700 228.9000 228.0700 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 109.9650 229.3400 230.4600 229.8400 ;
      RECT 108.5850 229.3400 109.4550 229.8400 ;
      RECT 107.2050 229.3400 108.0750 229.8400 ;
      RECT 105.8250 229.3400 106.6950 229.8400 ;
      RECT 104.4450 229.3400 105.3150 229.8400 ;
      RECT 103.0650 229.3400 103.9350 229.8400 ;
      RECT 101.6850 229.3400 102.5550 229.8400 ;
      RECT 100.3050 229.3400 101.1750 229.8400 ;
      RECT 98.9250 229.3400 99.7950 229.8400 ;
      RECT 98.0050 229.3400 98.4150 229.8400 ;
      RECT 96.6250 229.3400 97.4950 229.8400 ;
      RECT 95.2450 229.3400 96.1150 229.8400 ;
      RECT 93.8650 229.3400 94.7350 229.8400 ;
      RECT 92.4850 229.3400 93.3550 229.8400 ;
      RECT 91.1050 229.3400 91.9750 229.8400 ;
      RECT 89.7250 229.3400 90.5950 229.8400 ;
      RECT 88.3450 229.3400 89.2150 229.8400 ;
      RECT 86.9650 229.3400 87.8350 229.8400 ;
      RECT 86.0450 229.3400 86.4550 229.8400 ;
      RECT 84.6650 229.3400 85.5350 229.8400 ;
      RECT 83.2850 229.3400 84.1550 229.8400 ;
      RECT 81.9050 229.3400 82.7750 229.8400 ;
      RECT 80.5250 229.3400 81.3950 229.8400 ;
      RECT 79.1450 229.3400 80.0150 229.8400 ;
      RECT 77.7650 229.3400 78.6350 229.8400 ;
      RECT 76.3850 229.3400 77.2550 229.8400 ;
      RECT 75.0050 229.3400 75.8750 229.8400 ;
      RECT 74.0850 229.3400 74.4950 229.8400 ;
      RECT 72.7050 229.3400 73.5750 229.8400 ;
      RECT 71.3250 229.3400 72.1950 229.8400 ;
      RECT 69.9450 229.3400 70.8150 229.8400 ;
      RECT 68.5650 229.3400 69.4350 229.8400 ;
      RECT 67.1850 229.3400 68.0550 229.8400 ;
      RECT 65.8050 229.3400 66.6750 229.8400 ;
      RECT 64.4250 229.3400 65.2950 229.8400 ;
      RECT 63.0450 229.3400 63.9150 229.8400 ;
      RECT 62.1250 229.3400 62.5350 229.8400 ;
      RECT 60.7450 229.3400 61.6150 229.8400 ;
      RECT 59.3650 229.3400 60.2350 229.8400 ;
      RECT 57.9850 229.3400 58.8550 229.8400 ;
      RECT 56.6050 229.3400 57.4750 229.8400 ;
      RECT 55.2250 229.3400 56.0950 229.8400 ;
      RECT 53.8450 229.3400 54.7150 229.8400 ;
      RECT 52.4650 229.3400 53.3350 229.8400 ;
      RECT 51.0850 229.3400 51.9550 229.8400 ;
      RECT 50.1650 229.3400 50.5750 229.8400 ;
      RECT 48.7850 229.3400 49.6550 229.8400 ;
      RECT 47.4050 229.3400 48.2750 229.8400 ;
      RECT 46.0250 229.3400 46.8950 229.8400 ;
      RECT 44.6450 229.3400 45.5150 229.8400 ;
      RECT 43.2650 229.3400 44.1350 229.8400 ;
      RECT 41.8850 229.3400 42.7550 229.8400 ;
      RECT 40.5050 229.3400 41.3750 229.8400 ;
      RECT 39.1250 229.3400 39.9950 229.8400 ;
      RECT 38.2050 229.3400 38.6150 229.8400 ;
      RECT 36.8250 229.3400 37.6950 229.8400 ;
      RECT 35.4450 229.3400 36.3150 229.8400 ;
      RECT 34.0650 229.3400 34.9350 229.8400 ;
      RECT 32.6850 229.3400 33.5550 229.8400 ;
      RECT 31.3050 229.3400 32.1750 229.8400 ;
      RECT 29.9250 229.3400 30.7950 229.8400 ;
      RECT 28.5450 229.3400 29.4150 229.8400 ;
      RECT 27.1650 229.3400 28.0350 229.8400 ;
      RECT 26.2450 229.3400 26.6550 229.8400 ;
      RECT 24.8650 229.3400 25.7350 229.8400 ;
      RECT 23.4850 229.3400 24.3550 229.8400 ;
      RECT 22.1050 229.3400 22.9750 229.8400 ;
      RECT 20.7250 229.3400 21.5950 229.8400 ;
      RECT 19.3450 229.3400 20.2150 229.8400 ;
      RECT 17.9650 229.3400 18.8350 229.8400 ;
      RECT 16.5850 229.3400 17.4550 229.8400 ;
      RECT 15.6650 229.3400 16.0750 229.8400 ;
      RECT 0.0000 229.3400 15.1550 229.8400 ;
      RECT 0.0000 0.5000 230.4600 229.3400 ;
      RECT 109.9650 0.0000 230.4600 0.5000 ;
      RECT 108.5850 0.0000 109.4550 0.5000 ;
      RECT 107.2050 0.0000 108.0750 0.5000 ;
      RECT 105.8250 0.0000 106.6950 0.5000 ;
      RECT 104.4450 0.0000 105.3150 0.5000 ;
      RECT 103.0650 0.0000 103.9350 0.5000 ;
      RECT 101.6850 0.0000 102.5550 0.5000 ;
      RECT 100.3050 0.0000 101.1750 0.5000 ;
      RECT 98.9250 0.0000 99.7950 0.5000 ;
      RECT 98.0050 0.0000 98.4150 0.5000 ;
      RECT 96.6250 0.0000 97.4950 0.5000 ;
      RECT 95.2450 0.0000 96.1150 0.5000 ;
      RECT 93.8650 0.0000 94.7350 0.5000 ;
      RECT 92.4850 0.0000 93.3550 0.5000 ;
      RECT 91.1050 0.0000 91.9750 0.5000 ;
      RECT 89.7250 0.0000 90.5950 0.5000 ;
      RECT 88.3450 0.0000 89.2150 0.5000 ;
      RECT 86.9650 0.0000 87.8350 0.5000 ;
      RECT 86.0450 0.0000 86.4550 0.5000 ;
      RECT 84.6650 0.0000 85.5350 0.5000 ;
      RECT 83.2850 0.0000 84.1550 0.5000 ;
      RECT 81.9050 0.0000 82.7750 0.5000 ;
      RECT 80.5250 0.0000 81.3950 0.5000 ;
      RECT 79.1450 0.0000 80.0150 0.5000 ;
      RECT 77.7650 0.0000 78.6350 0.5000 ;
      RECT 76.3850 0.0000 77.2550 0.5000 ;
      RECT 75.0050 0.0000 75.8750 0.5000 ;
      RECT 74.0850 0.0000 74.4950 0.5000 ;
      RECT 72.7050 0.0000 73.5750 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 69.9450 0.0000 70.8150 0.5000 ;
      RECT 68.5650 0.0000 69.4350 0.5000 ;
      RECT 67.1850 0.0000 68.0550 0.5000 ;
      RECT 65.8050 0.0000 66.6750 0.5000 ;
      RECT 64.4250 0.0000 65.2950 0.5000 ;
      RECT 63.0450 0.0000 63.9150 0.5000 ;
      RECT 62.1250 0.0000 62.5350 0.5000 ;
      RECT 60.7450 0.0000 61.6150 0.5000 ;
      RECT 59.3650 0.0000 60.2350 0.5000 ;
      RECT 57.9850 0.0000 58.8550 0.5000 ;
      RECT 56.6050 0.0000 57.4750 0.5000 ;
      RECT 55.2250 0.0000 56.0950 0.5000 ;
      RECT 53.8450 0.0000 54.7150 0.5000 ;
      RECT 52.4650 0.0000 53.3350 0.5000 ;
      RECT 51.0850 0.0000 51.9550 0.5000 ;
      RECT 50.1650 0.0000 50.5750 0.5000 ;
      RECT 48.7850 0.0000 49.6550 0.5000 ;
      RECT 47.4050 0.0000 48.2750 0.5000 ;
      RECT 46.0250 0.0000 46.8950 0.5000 ;
      RECT 44.6450 0.0000 45.5150 0.5000 ;
      RECT 43.2650 0.0000 44.1350 0.5000 ;
      RECT 41.8850 0.0000 42.7550 0.5000 ;
      RECT 40.5050 0.0000 41.3750 0.5000 ;
      RECT 39.1250 0.0000 39.9950 0.5000 ;
      RECT 38.2050 0.0000 38.6150 0.5000 ;
      RECT 36.8250 0.0000 37.6950 0.5000 ;
      RECT 35.4450 0.0000 36.3150 0.5000 ;
      RECT 34.0650 0.0000 34.9350 0.5000 ;
      RECT 32.6850 0.0000 33.5550 0.5000 ;
      RECT 31.3050 0.0000 32.1750 0.5000 ;
      RECT 29.9250 0.0000 30.7950 0.5000 ;
      RECT 28.5450 0.0000 29.4150 0.5000 ;
      RECT 27.1650 0.0000 28.0350 0.5000 ;
      RECT 26.2450 0.0000 26.6550 0.5000 ;
      RECT 24.8650 0.0000 25.7350 0.5000 ;
      RECT 23.4850 0.0000 24.3550 0.5000 ;
      RECT 22.1050 0.0000 22.9750 0.5000 ;
      RECT 20.7250 0.0000 21.5950 0.5000 ;
      RECT 19.3450 0.0000 20.2150 0.5000 ;
      RECT 17.9650 0.0000 18.8350 0.5000 ;
      RECT 16.5850 0.0000 17.4550 0.5000 ;
      RECT 15.6650 0.0000 16.0750 0.5000 ;
      RECT 0.0000 0.0000 15.1550 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 230.4600 229.8400 ;
    LAYER met2 ;
      RECT 214.8000 229.2150 230.4600 229.8400 ;
      RECT 209.2800 229.2150 214.3800 229.8400 ;
      RECT 205.1400 229.2150 208.8600 229.8400 ;
      RECT 200.5400 229.2150 204.7200 229.8400 ;
      RECT 195.9400 229.2150 200.1200 229.8400 ;
      RECT 190.8800 229.2150 195.5200 229.8400 ;
      RECT 186.2800 229.2150 190.4600 229.8400 ;
      RECT 181.6800 229.2150 185.8600 229.8400 ;
      RECT 177.0800 229.2150 181.2600 229.8400 ;
      RECT 172.0200 229.2150 176.6600 229.8400 ;
      RECT 167.4200 229.2150 171.6000 229.8400 ;
      RECT 162.8200 229.2150 167.0000 229.8400 ;
      RECT 158.2200 229.2150 162.4000 229.8400 ;
      RECT 153.1600 229.2150 157.8000 229.8400 ;
      RECT 148.5600 229.2150 152.7400 229.8400 ;
      RECT 143.9600 229.2150 148.1400 229.8400 ;
      RECT 139.3600 229.2150 143.5400 229.8400 ;
      RECT 134.3000 229.2150 138.9400 229.8400 ;
      RECT 129.7000 229.2150 133.8800 229.8400 ;
      RECT 125.1000 229.2150 129.2800 229.8400 ;
      RECT 120.5000 229.2150 124.6800 229.8400 ;
      RECT 0.0000 229.2150 120.0800 229.8400 ;
      RECT 0.0000 228.2100 230.4600 229.2150 ;
      RECT 195.0600 224.2100 225.7600 228.2100 ;
      RECT 165.0600 224.2100 193.1800 228.2100 ;
      RECT 135.0600 224.2100 163.1800 228.2100 ;
      RECT 105.0600 224.2100 133.1800 228.2100 ;
      RECT 75.0600 224.2100 103.1800 228.2100 ;
      RECT 45.0600 224.2100 73.1800 228.2100 ;
      RECT 15.0600 224.2100 43.1800 228.2100 ;
      RECT 4.7000 224.2100 13.1800 228.2100 ;
      RECT 229.0400 214.5800 230.4600 228.2100 ;
      RECT 0.0000 214.5800 1.4200 228.2100 ;
      RECT 229.0400 214.1600 229.8350 214.5800 ;
      RECT 0.6250 214.1600 1.4200 214.5800 ;
      RECT 229.0400 211.8600 230.4600 214.1600 ;
      RECT 0.0000 211.8600 1.4200 214.1600 ;
      RECT 229.0400 211.4400 229.8350 211.8600 ;
      RECT 0.6250 211.4400 1.4200 211.8600 ;
      RECT 229.0400 208.8000 230.4600 211.4400 ;
      RECT 0.0000 208.8000 1.4200 211.4400 ;
      RECT 229.0400 208.3800 229.8350 208.8000 ;
      RECT 0.6250 208.3800 1.4200 208.8000 ;
      RECT 229.0400 205.7400 230.4600 208.3800 ;
      RECT 0.0000 205.7400 1.4200 208.3800 ;
      RECT 229.0400 205.3200 229.8350 205.7400 ;
      RECT 0.6250 205.3200 1.4200 205.7400 ;
      RECT 229.0400 202.6800 230.4600 205.3200 ;
      RECT 0.0000 202.6800 1.4200 205.3200 ;
      RECT 229.0400 202.2600 229.8350 202.6800 ;
      RECT 0.6250 202.2600 1.4200 202.6800 ;
      RECT 229.0400 199.6200 230.4600 202.2600 ;
      RECT 0.0000 199.6200 1.4200 202.2600 ;
      RECT 229.0400 199.2000 229.8350 199.6200 ;
      RECT 0.6250 199.2000 1.4200 199.6200 ;
      RECT 229.0400 196.5600 230.4600 199.2000 ;
      RECT 0.0000 196.5600 1.4200 199.2000 ;
      RECT 229.0400 196.1400 229.8350 196.5600 ;
      RECT 0.6250 196.1400 1.4200 196.5600 ;
      RECT 229.0400 193.5000 230.4600 196.1400 ;
      RECT 0.0000 193.5000 1.4200 196.1400 ;
      RECT 229.0400 193.0800 229.8350 193.5000 ;
      RECT 0.6250 193.0800 1.4200 193.5000 ;
      RECT 229.0400 190.4400 230.4600 193.0800 ;
      RECT 0.0000 190.4400 1.4200 193.0800 ;
      RECT 229.0400 190.0200 229.8350 190.4400 ;
      RECT 0.6250 190.0200 1.4200 190.4400 ;
      RECT 229.0400 187.3800 230.4600 190.0200 ;
      RECT 0.0000 187.3800 1.4200 190.0200 ;
      RECT 229.0400 186.9600 229.8350 187.3800 ;
      RECT 0.6250 186.9600 1.4200 187.3800 ;
      RECT 229.0400 184.3200 230.4600 186.9600 ;
      RECT 0.0000 184.3200 1.4200 186.9600 ;
      RECT 229.0400 183.9000 229.8350 184.3200 ;
      RECT 0.6250 183.9000 1.4200 184.3200 ;
      RECT 229.0400 181.2600 230.4600 183.9000 ;
      RECT 0.0000 181.2600 1.4200 183.9000 ;
      RECT 229.0400 180.8400 229.8350 181.2600 ;
      RECT 0.6250 180.8400 1.4200 181.2600 ;
      RECT 229.0400 178.2000 230.4600 180.8400 ;
      RECT 0.0000 178.2000 1.4200 180.8400 ;
      RECT 229.0400 177.7800 229.8350 178.2000 ;
      RECT 0.6250 177.7800 1.4200 178.2000 ;
      RECT 229.0400 175.1400 230.4600 177.7800 ;
      RECT 0.0000 175.1400 1.4200 177.7800 ;
      RECT 229.0400 174.7200 229.8350 175.1400 ;
      RECT 0.6250 174.7200 1.4200 175.1400 ;
      RECT 229.0400 172.0800 230.4600 174.7200 ;
      RECT 0.0000 172.0800 1.4200 174.7200 ;
      RECT 229.0400 171.6600 229.8350 172.0800 ;
      RECT 0.6250 171.6600 1.4200 172.0800 ;
      RECT 229.0400 169.0200 230.4600 171.6600 ;
      RECT 0.0000 169.0200 1.4200 171.6600 ;
      RECT 229.0400 168.6000 229.8350 169.0200 ;
      RECT 0.6250 168.6000 1.4200 169.0200 ;
      RECT 229.0400 165.9600 230.4600 168.6000 ;
      RECT 0.0000 165.9600 1.4200 168.6000 ;
      RECT 229.0400 165.5400 229.8350 165.9600 ;
      RECT 0.6250 165.5400 1.4200 165.9600 ;
      RECT 229.0400 162.9000 230.4600 165.5400 ;
      RECT 0.0000 162.9000 1.4200 165.5400 ;
      RECT 229.0400 162.4800 229.8350 162.9000 ;
      RECT 0.6250 162.4800 1.4200 162.9000 ;
      RECT 229.0400 159.8400 230.4600 162.4800 ;
      RECT 0.0000 159.8400 1.4200 162.4800 ;
      RECT 229.0400 159.4200 229.8350 159.8400 ;
      RECT 0.6250 159.4200 1.4200 159.8400 ;
      RECT 229.0400 156.7800 230.4600 159.4200 ;
      RECT 0.0000 156.7800 1.4200 159.4200 ;
      RECT 229.0400 156.3600 229.8350 156.7800 ;
      RECT 0.6250 156.3600 1.4200 156.7800 ;
      RECT 229.0400 153.7200 230.4600 156.3600 ;
      RECT 0.0000 153.7200 1.4200 156.3600 ;
      RECT 229.0400 153.3000 229.8350 153.7200 ;
      RECT 0.6250 153.3000 1.4200 153.7200 ;
      RECT 229.0400 150.6600 230.4600 153.3000 ;
      RECT 0.0000 150.6600 1.4200 153.3000 ;
      RECT 229.0400 150.2400 229.8350 150.6600 ;
      RECT 0.6250 150.2400 1.4200 150.6600 ;
      RECT 229.0400 147.6000 230.4600 150.2400 ;
      RECT 0.0000 147.6000 1.4200 150.2400 ;
      RECT 229.0400 147.1800 229.8350 147.6000 ;
      RECT 0.6250 147.1800 1.4200 147.6000 ;
      RECT 229.0400 144.5400 230.4600 147.1800 ;
      RECT 0.0000 144.5400 1.4200 147.1800 ;
      RECT 229.0400 144.1200 229.8350 144.5400 ;
      RECT 0.6250 144.1200 1.4200 144.5400 ;
      RECT 229.0400 141.4800 230.4600 144.1200 ;
      RECT 0.0000 141.4800 1.4200 144.1200 ;
      RECT 229.0400 141.0600 229.8350 141.4800 ;
      RECT 0.6250 141.0600 1.4200 141.4800 ;
      RECT 229.0400 138.4200 230.4600 141.0600 ;
      RECT 0.0000 138.4200 1.4200 141.0600 ;
      RECT 229.0400 138.0000 229.8350 138.4200 ;
      RECT 0.6250 138.0000 1.4200 138.4200 ;
      RECT 229.0400 135.3600 230.4600 138.0000 ;
      RECT 0.0000 135.3600 1.4200 138.0000 ;
      RECT 229.0400 134.9400 229.8350 135.3600 ;
      RECT 0.6250 134.9400 1.4200 135.3600 ;
      RECT 229.0400 132.3000 230.4600 134.9400 ;
      RECT 0.0000 132.3000 1.4200 134.9400 ;
      RECT 229.0400 131.8800 229.8350 132.3000 ;
      RECT 0.6250 131.8800 1.4200 132.3000 ;
      RECT 229.0400 129.2400 230.4600 131.8800 ;
      RECT 0.0000 129.2400 1.4200 131.8800 ;
      RECT 229.0400 128.8200 229.8350 129.2400 ;
      RECT 0.6250 128.8200 1.4200 129.2400 ;
      RECT 229.0400 126.1800 230.4600 128.8200 ;
      RECT 0.0000 126.1800 1.4200 128.8200 ;
      RECT 229.0400 125.7600 229.8350 126.1800 ;
      RECT 0.6250 125.7600 1.4200 126.1800 ;
      RECT 229.0400 123.1200 230.4600 125.7600 ;
      RECT 0.0000 123.1200 1.4200 125.7600 ;
      RECT 229.0400 122.7000 229.8350 123.1200 ;
      RECT 0.6250 122.7000 1.4200 123.1200 ;
      RECT 229.0400 120.4000 230.4600 122.7000 ;
      RECT 0.0000 120.4000 1.4200 122.7000 ;
      RECT 229.0400 119.9800 229.8350 120.4000 ;
      RECT 0.6250 119.9800 1.4200 120.4000 ;
      RECT 229.0400 109.8600 230.4600 119.9800 ;
      RECT 0.0000 109.8600 1.4200 119.9800 ;
      RECT 229.0400 109.4400 229.8350 109.8600 ;
      RECT 0.6250 109.4400 1.4200 109.8600 ;
      RECT 229.0400 108.5000 230.4600 109.4400 ;
      RECT 0.0000 108.5000 1.4200 109.4400 ;
      RECT 229.0400 108.0800 229.8350 108.5000 ;
      RECT 0.6250 108.0800 1.4200 108.5000 ;
      RECT 229.0400 107.1400 230.4600 108.0800 ;
      RECT 0.0000 107.1400 1.4200 108.0800 ;
      RECT 229.0400 106.7200 229.8350 107.1400 ;
      RECT 0.6250 106.7200 1.4200 107.1400 ;
      RECT 229.0400 105.4400 230.4600 106.7200 ;
      RECT 0.0000 105.4400 1.4200 106.7200 ;
      RECT 229.0400 105.0200 229.8350 105.4400 ;
      RECT 0.6250 105.0200 1.4200 105.4400 ;
      RECT 229.0400 104.0800 230.4600 105.0200 ;
      RECT 0.0000 104.0800 1.4200 105.0200 ;
      RECT 229.0400 103.6600 229.8350 104.0800 ;
      RECT 0.6250 103.6600 1.4200 104.0800 ;
      RECT 229.0400 102.3800 230.4600 103.6600 ;
      RECT 0.0000 102.3800 1.4200 103.6600 ;
      RECT 229.0400 101.9600 229.8350 102.3800 ;
      RECT 0.6250 101.9600 1.4200 102.3800 ;
      RECT 229.0400 101.0200 230.4600 101.9600 ;
      RECT 0.0000 101.0200 1.4200 101.9600 ;
      RECT 229.0400 100.6000 229.8350 101.0200 ;
      RECT 0.6250 100.6000 1.4200 101.0200 ;
      RECT 229.0400 99.3200 230.4600 100.6000 ;
      RECT 0.0000 99.3200 1.4200 100.6000 ;
      RECT 229.0400 98.9000 229.8350 99.3200 ;
      RECT 0.6250 98.9000 1.4200 99.3200 ;
      RECT 229.0400 97.9600 230.4600 98.9000 ;
      RECT 0.0000 97.9600 1.4200 98.9000 ;
      RECT 229.0400 97.5400 229.8350 97.9600 ;
      RECT 0.6250 97.5400 1.4200 97.9600 ;
      RECT 229.0400 96.6000 230.4600 97.5400 ;
      RECT 0.0000 96.6000 1.4200 97.5400 ;
      RECT 229.0400 96.1800 229.8350 96.6000 ;
      RECT 0.6250 96.1800 1.4200 96.6000 ;
      RECT 229.0400 94.9000 230.4600 96.1800 ;
      RECT 0.0000 94.9000 1.4200 96.1800 ;
      RECT 229.0400 94.4800 229.8350 94.9000 ;
      RECT 0.6250 94.4800 1.4200 94.9000 ;
      RECT 229.0400 93.5400 230.4600 94.4800 ;
      RECT 0.0000 93.5400 1.4200 94.4800 ;
      RECT 229.0400 93.1200 229.8350 93.5400 ;
      RECT 0.6250 93.1200 1.4200 93.5400 ;
      RECT 229.0400 91.8400 230.4600 93.1200 ;
      RECT 0.0000 91.8400 1.4200 93.1200 ;
      RECT 229.0400 91.4200 229.8350 91.8400 ;
      RECT 0.6250 91.4200 1.4200 91.8400 ;
      RECT 229.0400 90.4800 230.4600 91.4200 ;
      RECT 0.0000 90.4800 1.4200 91.4200 ;
      RECT 229.0400 90.0600 229.8350 90.4800 ;
      RECT 0.6250 90.0600 1.4200 90.4800 ;
      RECT 229.0400 88.7800 230.4600 90.0600 ;
      RECT 0.0000 88.7800 1.4200 90.0600 ;
      RECT 229.0400 88.3600 229.8350 88.7800 ;
      RECT 0.6250 88.3600 1.4200 88.7800 ;
      RECT 229.0400 87.4200 230.4600 88.3600 ;
      RECT 0.0000 87.4200 1.4200 88.3600 ;
      RECT 229.0400 87.0000 229.8350 87.4200 ;
      RECT 0.6250 87.0000 1.4200 87.4200 ;
      RECT 229.0400 86.0600 230.4600 87.0000 ;
      RECT 0.0000 86.0600 1.4200 87.0000 ;
      RECT 229.0400 85.6400 229.8350 86.0600 ;
      RECT 0.6250 85.6400 1.4200 86.0600 ;
      RECT 229.0400 84.3600 230.4600 85.6400 ;
      RECT 0.0000 84.3600 1.4200 85.6400 ;
      RECT 229.0400 83.9400 229.8350 84.3600 ;
      RECT 0.6250 83.9400 1.4200 84.3600 ;
      RECT 229.0400 83.0000 230.4600 83.9400 ;
      RECT 0.0000 83.0000 1.4200 83.9400 ;
      RECT 229.0400 82.5800 229.8350 83.0000 ;
      RECT 0.6250 82.5800 1.4200 83.0000 ;
      RECT 229.0400 81.3000 230.4600 82.5800 ;
      RECT 0.0000 81.3000 1.4200 82.5800 ;
      RECT 229.0400 80.8800 229.8350 81.3000 ;
      RECT 0.6250 80.8800 1.4200 81.3000 ;
      RECT 229.0400 79.9400 230.4600 80.8800 ;
      RECT 0.0000 79.9400 1.4200 80.8800 ;
      RECT 229.0400 79.5200 229.8350 79.9400 ;
      RECT 0.6250 79.5200 1.4200 79.9400 ;
      RECT 229.0400 78.2400 230.4600 79.5200 ;
      RECT 0.0000 78.2400 1.4200 79.5200 ;
      RECT 229.0400 77.8200 229.8350 78.2400 ;
      RECT 0.6250 77.8200 1.4200 78.2400 ;
      RECT 229.0400 76.8800 230.4600 77.8200 ;
      RECT 0.0000 76.8800 1.4200 77.8200 ;
      RECT 229.0400 76.4600 229.8350 76.8800 ;
      RECT 0.6250 76.4600 1.4200 76.8800 ;
      RECT 229.0400 75.5200 230.4600 76.4600 ;
      RECT 0.0000 75.5200 1.4200 76.4600 ;
      RECT 229.0400 75.1000 229.8350 75.5200 ;
      RECT 0.6250 75.1000 1.4200 75.5200 ;
      RECT 229.0400 73.8200 230.4600 75.1000 ;
      RECT 0.0000 73.8200 1.4200 75.1000 ;
      RECT 229.0400 73.4000 229.8350 73.8200 ;
      RECT 0.6250 73.4000 1.4200 73.8200 ;
      RECT 229.0400 72.4600 230.4600 73.4000 ;
      RECT 0.0000 72.4600 1.4200 73.4000 ;
      RECT 229.0400 72.0400 229.8350 72.4600 ;
      RECT 0.6250 72.0400 1.4200 72.4600 ;
      RECT 229.0400 70.7600 230.4600 72.0400 ;
      RECT 0.0000 70.7600 1.4200 72.0400 ;
      RECT 229.0400 70.3400 229.8350 70.7600 ;
      RECT 0.6250 70.3400 1.4200 70.7600 ;
      RECT 229.0400 69.4000 230.4600 70.3400 ;
      RECT 0.0000 69.4000 1.4200 70.3400 ;
      RECT 229.0400 68.9800 229.8350 69.4000 ;
      RECT 0.6250 68.9800 1.4200 69.4000 ;
      RECT 229.0400 67.7000 230.4600 68.9800 ;
      RECT 0.0000 67.7000 1.4200 68.9800 ;
      RECT 229.0400 67.2800 229.8350 67.7000 ;
      RECT 0.6250 67.2800 1.4200 67.7000 ;
      RECT 229.0400 66.3400 230.4600 67.2800 ;
      RECT 0.0000 66.3400 1.4200 67.2800 ;
      RECT 229.0400 65.9200 229.8350 66.3400 ;
      RECT 0.6250 65.9200 1.4200 66.3400 ;
      RECT 229.0400 64.9800 230.4600 65.9200 ;
      RECT 0.0000 64.9800 1.4200 65.9200 ;
      RECT 229.0400 64.5600 229.8350 64.9800 ;
      RECT 0.6250 64.5600 1.4200 64.9800 ;
      RECT 229.0400 63.2800 230.4600 64.5600 ;
      RECT 0.0000 63.2800 1.4200 64.5600 ;
      RECT 229.0400 62.8600 229.8350 63.2800 ;
      RECT 0.6250 62.8600 1.4200 63.2800 ;
      RECT 229.0400 61.9200 230.4600 62.8600 ;
      RECT 0.0000 61.9200 1.4200 62.8600 ;
      RECT 229.0400 61.5000 229.8350 61.9200 ;
      RECT 0.6250 61.5000 1.4200 61.9200 ;
      RECT 229.0400 60.2200 230.4600 61.5000 ;
      RECT 0.0000 60.2200 1.4200 61.5000 ;
      RECT 229.0400 59.8000 229.8350 60.2200 ;
      RECT 0.6250 59.8000 1.4200 60.2200 ;
      RECT 229.0400 58.8600 230.4600 59.8000 ;
      RECT 0.0000 58.8600 1.4200 59.8000 ;
      RECT 229.0400 58.4400 229.8350 58.8600 ;
      RECT 0.6250 58.4400 1.4200 58.8600 ;
      RECT 229.0400 57.5000 230.4600 58.4400 ;
      RECT 0.0000 57.5000 1.4200 58.4400 ;
      RECT 229.0400 57.0800 229.8350 57.5000 ;
      RECT 0.6250 57.0800 1.4200 57.5000 ;
      RECT 229.0400 55.8000 230.4600 57.0800 ;
      RECT 0.0000 55.8000 1.4200 57.0800 ;
      RECT 229.0400 55.3800 229.8350 55.8000 ;
      RECT 0.6250 55.3800 1.4200 55.8000 ;
      RECT 229.0400 54.4400 230.4600 55.3800 ;
      RECT 0.0000 54.4400 1.4200 55.3800 ;
      RECT 229.0400 54.0200 229.8350 54.4400 ;
      RECT 0.6250 54.0200 1.4200 54.4400 ;
      RECT 229.0400 52.7400 230.4600 54.0200 ;
      RECT 0.0000 52.7400 1.4200 54.0200 ;
      RECT 229.0400 52.3200 229.8350 52.7400 ;
      RECT 0.6250 52.3200 1.4200 52.7400 ;
      RECT 229.0400 51.3800 230.4600 52.3200 ;
      RECT 0.0000 51.3800 1.4200 52.3200 ;
      RECT 229.0400 50.9600 229.8350 51.3800 ;
      RECT 0.6250 50.9600 1.4200 51.3800 ;
      RECT 229.0400 49.6800 230.4600 50.9600 ;
      RECT 0.0000 49.6800 1.4200 50.9600 ;
      RECT 229.0400 49.2600 229.8350 49.6800 ;
      RECT 0.6250 49.2600 1.4200 49.6800 ;
      RECT 229.0400 48.3200 230.4600 49.2600 ;
      RECT 0.0000 48.3200 1.4200 49.2600 ;
      RECT 229.0400 47.9000 229.8350 48.3200 ;
      RECT 0.6250 47.9000 1.4200 48.3200 ;
      RECT 229.0400 46.9600 230.4600 47.9000 ;
      RECT 0.0000 46.9600 1.4200 47.9000 ;
      RECT 229.0400 46.5400 229.8350 46.9600 ;
      RECT 0.6250 46.5400 1.4200 46.9600 ;
      RECT 229.0400 45.2600 230.4600 46.5400 ;
      RECT 0.0000 45.2600 1.4200 46.5400 ;
      RECT 229.0400 44.8400 229.8350 45.2600 ;
      RECT 0.6250 44.8400 1.4200 45.2600 ;
      RECT 229.0400 43.9000 230.4600 44.8400 ;
      RECT 0.0000 43.9000 1.4200 44.8400 ;
      RECT 229.0400 43.4800 229.8350 43.9000 ;
      RECT 0.6250 43.4800 1.4200 43.9000 ;
      RECT 229.0400 42.2000 230.4600 43.4800 ;
      RECT 0.0000 42.2000 1.4200 43.4800 ;
      RECT 229.0400 41.7800 229.8350 42.2000 ;
      RECT 0.6250 41.7800 1.4200 42.2000 ;
      RECT 229.0400 40.8400 230.4600 41.7800 ;
      RECT 0.0000 40.8400 1.4200 41.7800 ;
      RECT 229.0400 40.4200 229.8350 40.8400 ;
      RECT 0.6250 40.4200 1.4200 40.8400 ;
      RECT 229.0400 39.1400 230.4600 40.4200 ;
      RECT 0.0000 39.1400 1.4200 40.4200 ;
      RECT 229.0400 38.7200 229.8350 39.1400 ;
      RECT 0.6250 38.7200 1.4200 39.1400 ;
      RECT 229.0400 37.7800 230.4600 38.7200 ;
      RECT 0.0000 37.7800 1.4200 38.7200 ;
      RECT 229.0400 37.3600 229.8350 37.7800 ;
      RECT 0.6250 37.3600 1.4200 37.7800 ;
      RECT 229.0400 36.4200 230.4600 37.3600 ;
      RECT 0.0000 36.4200 1.4200 37.3600 ;
      RECT 229.0400 36.0000 229.8350 36.4200 ;
      RECT 0.6250 36.0000 1.4200 36.4200 ;
      RECT 229.0400 34.7200 230.4600 36.0000 ;
      RECT 0.0000 34.7200 1.4200 36.0000 ;
      RECT 229.0400 34.3000 229.8350 34.7200 ;
      RECT 0.6250 34.3000 1.4200 34.7200 ;
      RECT 229.0400 33.3600 230.4600 34.3000 ;
      RECT 0.0000 33.3600 1.4200 34.3000 ;
      RECT 229.0400 32.9400 229.8350 33.3600 ;
      RECT 0.6250 32.9400 1.4200 33.3600 ;
      RECT 229.0400 31.6600 230.4600 32.9400 ;
      RECT 0.0000 31.6600 1.4200 32.9400 ;
      RECT 229.0400 31.2400 229.8350 31.6600 ;
      RECT 0.6250 31.2400 1.4200 31.6600 ;
      RECT 229.0400 30.3000 230.4600 31.2400 ;
      RECT 0.0000 30.3000 1.4200 31.2400 ;
      RECT 229.0400 29.8800 229.8350 30.3000 ;
      RECT 0.6250 29.8800 1.4200 30.3000 ;
      RECT 229.0400 28.6000 230.4600 29.8800 ;
      RECT 0.0000 28.6000 1.4200 29.8800 ;
      RECT 229.0400 28.1800 229.8350 28.6000 ;
      RECT 0.6250 28.1800 1.4200 28.6000 ;
      RECT 229.0400 27.2400 230.4600 28.1800 ;
      RECT 0.0000 27.2400 1.4200 28.1800 ;
      RECT 229.0400 26.8200 229.8350 27.2400 ;
      RECT 0.6250 26.8200 1.4200 27.2400 ;
      RECT 229.0400 25.8800 230.4600 26.8200 ;
      RECT 0.0000 25.8800 1.4200 26.8200 ;
      RECT 229.0400 25.4600 229.8350 25.8800 ;
      RECT 0.6250 25.4600 1.4200 25.8800 ;
      RECT 229.0400 24.1800 230.4600 25.4600 ;
      RECT 0.0000 24.1800 1.4200 25.4600 ;
      RECT 229.0400 23.7600 229.8350 24.1800 ;
      RECT 0.6250 23.7600 1.4200 24.1800 ;
      RECT 229.0400 22.8200 230.4600 23.7600 ;
      RECT 0.0000 22.8200 1.4200 23.7600 ;
      RECT 229.0400 22.4000 229.8350 22.8200 ;
      RECT 0.6250 22.4000 1.4200 22.8200 ;
      RECT 229.0400 21.1200 230.4600 22.4000 ;
      RECT 0.0000 21.1200 1.4200 22.4000 ;
      RECT 229.0400 20.7000 229.8350 21.1200 ;
      RECT 0.6250 20.7000 1.4200 21.1200 ;
      RECT 229.0400 19.7600 230.4600 20.7000 ;
      RECT 0.0000 19.7600 1.4200 20.7000 ;
      RECT 229.0400 19.3400 229.8350 19.7600 ;
      RECT 0.6250 19.3400 1.4200 19.7600 ;
      RECT 229.0400 18.0600 230.4600 19.3400 ;
      RECT 0.0000 18.0600 1.4200 19.3400 ;
      RECT 229.0400 17.6400 229.8350 18.0600 ;
      RECT 0.6250 17.6400 1.4200 18.0600 ;
      RECT 229.0400 16.7000 230.4600 17.6400 ;
      RECT 0.0000 16.7000 1.4200 17.6400 ;
      RECT 229.0400 16.2800 229.8350 16.7000 ;
      RECT 0.6250 16.2800 1.4200 16.7000 ;
      RECT 229.0400 15.3400 230.4600 16.2800 ;
      RECT 0.0000 15.3400 1.4200 16.2800 ;
      RECT 229.0400 14.9200 229.8350 15.3400 ;
      RECT 0.6250 14.9200 1.4200 15.3400 ;
      RECT 225.0400 5.2900 225.7600 224.2100 ;
      RECT 195.0600 5.2900 221.7600 224.2100 ;
      RECT 191.8600 5.2900 193.1800 224.2100 ;
      RECT 165.0600 5.2900 189.9800 224.2100 ;
      RECT 161.8600 5.2900 163.1800 224.2100 ;
      RECT 135.0600 5.2900 159.9800 224.2100 ;
      RECT 131.8600 5.2900 133.1800 224.2100 ;
      RECT 105.0600 5.2900 129.9800 224.2100 ;
      RECT 101.8600 5.2900 103.1800 224.2100 ;
      RECT 75.0600 5.2900 99.9800 224.2100 ;
      RECT 71.8600 5.2900 73.1800 224.2100 ;
      RECT 45.0600 5.2900 69.9800 224.2100 ;
      RECT 41.8600 5.2900 43.1800 224.2100 ;
      RECT 15.0600 5.2900 39.9800 224.2100 ;
      RECT 8.7000 5.2900 13.1800 224.2100 ;
      RECT 4.7000 5.2900 5.4200 224.2100 ;
      RECT 229.0400 1.2900 230.4600 14.9200 ;
      RECT 195.0600 1.2900 225.7600 5.2900 ;
      RECT 165.0600 1.2900 193.1800 5.2900 ;
      RECT 135.0600 1.2900 163.1800 5.2900 ;
      RECT 105.0600 1.2900 133.1800 5.2900 ;
      RECT 75.0600 1.2900 103.1800 5.2900 ;
      RECT 45.0600 1.2900 73.1800 5.2900 ;
      RECT 15.0600 1.2900 43.1800 5.2900 ;
      RECT 4.7000 1.2900 13.1800 5.2900 ;
      RECT 0.0000 1.2900 1.4200 14.9200 ;
      RECT 0.0000 0.6250 230.4600 1.2900 ;
      RECT 214.3400 0.0000 230.4600 0.6250 ;
      RECT 209.7400 0.0000 213.9200 0.6250 ;
      RECT 205.1400 0.0000 209.3200 0.6250 ;
      RECT 200.5400 0.0000 204.7200 0.6250 ;
      RECT 195.9400 0.0000 200.1200 0.6250 ;
      RECT 191.3400 0.0000 195.5200 0.6250 ;
      RECT 186.2800 0.0000 190.9200 0.6250 ;
      RECT 181.6800 0.0000 185.8600 0.6250 ;
      RECT 177.0800 0.0000 181.2600 0.6250 ;
      RECT 172.4800 0.0000 176.6600 0.6250 ;
      RECT 167.8800 0.0000 172.0600 0.6250 ;
      RECT 162.8200 0.0000 167.4600 0.6250 ;
      RECT 158.2200 0.0000 162.4000 0.6250 ;
      RECT 153.6200 0.0000 157.8000 0.6250 ;
      RECT 149.0200 0.0000 153.2000 0.6250 ;
      RECT 144.4200 0.0000 148.6000 0.6250 ;
      RECT 139.3600 0.0000 144.0000 0.6250 ;
      RECT 134.7600 0.0000 138.9400 0.6250 ;
      RECT 129.7000 0.0000 134.3400 0.6250 ;
      RECT 125.5600 0.0000 129.2800 0.6250 ;
      RECT 120.9600 0.0000 125.1400 0.6250 ;
      RECT 0.0000 0.0000 120.5400 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 228.3700 230.4600 229.8400 ;
      RECT 229.2000 224.7700 230.4600 228.3700 ;
      RECT 0.0000 224.7700 1.2600 228.3700 ;
      RECT 0.0000 224.3700 230.4600 224.7700 ;
      RECT 225.2000 220.7700 230.4600 224.3700 ;
      RECT 0.0000 220.7700 5.2600 224.3700 ;
      RECT 0.0000 8.7300 230.4600 220.7700 ;
      RECT 225.2000 5.1300 230.4600 8.7300 ;
      RECT 0.0000 5.1300 5.2600 8.7300 ;
      RECT 0.0000 4.7300 230.4600 5.1300 ;
      RECT 229.2000 1.1300 230.4600 4.7300 ;
      RECT 0.0000 1.1300 1.2600 4.7300 ;
      RECT 0.0000 0.0000 230.4600 1.1300 ;
  END
END LUT4AB

END LIBRARY
