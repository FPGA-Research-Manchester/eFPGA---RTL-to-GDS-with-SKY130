##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Wed Apr 21 17:46:52 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO W_IO
  CLASS BLOCK ;
  SIZE 29.9000 BY 229.8400 ;
  FOREIGN W_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5533 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6215 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.1166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.347 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 67.4200 29.9000 67.5600 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8777 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.808 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 66.0600 29.9000 66.2000 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6729 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.662 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 64.7000 29.9000 64.8400 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.2418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.76 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 63.0000 29.9000 63.1400 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.0681 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.236 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 79.6600 29.9000 79.8000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.0397 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.131 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 77.9600 29.9000 78.1000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7657 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 76.6000 29.9000 76.7400 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.9592 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7285 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 75.2400 29.9000 75.3800 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3285 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.896 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 73.5400 29.9000 73.6800 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4405 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.3556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.66 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 72.1800 29.9000 72.3200 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.4856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.31 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 70.4800 29.9000 70.6200 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.9795 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.83 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 69.1200 29.9000 69.2600 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.0068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 91.5600 29.9000 91.7000 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.0415 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.103 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 90.2000 29.9000 90.3400 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.9897 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.844 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 88.5000 29.9000 88.6400 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.9277 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.571 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 87.1400 29.9000 87.2800 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.116 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.66 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 85.7800 29.9000 85.9200 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.53 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 84.0800 29.9000 84.2200 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.7681 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.773 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 82.7200 29.9000 82.8600 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 0.9897 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.844 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 81.0200 29.9000 81.1600 ;
    END
  END E2BEGb[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7097 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4035 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.076 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 109.5800 29.9000 109.7200 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.61 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.152 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 108.2200 29.9000 108.3600 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.9095 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 106.8600 29.9000 107.0000 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0993 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3515 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.054 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 105.1600 29.9000 105.3000 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.8619 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.205 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 103.8000 29.9000 103.9400 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.262 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.1184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.474 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 102.1000 29.9000 102.2400 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.1157 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.474 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 100.7400 29.9000 100.8800 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.284 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 99.0400 29.9000 99.1800 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 97.6800 29.9000 97.8200 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3401 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 96.3200 29.9000 96.4600 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3779 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 94.6200 29.9000 94.7600 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.1543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.6005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 3.564 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.8938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 93.2600 29.9000 93.4000 ;
    END
  END E6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 19.4800 29.9000 19.6200 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 17.7800 29.9000 17.9200 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 16.4200 29.9000 16.5600 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 15.0600 29.9000 15.2000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2112 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.948 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.9652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.482 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.98 LAYER met2  ;
    ANTENNAMAXAREACAR 5.54848 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.9859 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 31.3800 29.9000 31.5200 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.1968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.98 LAYER met4  ;
    ANTENNAMAXAREACAR 36.5371 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 183.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.64202 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 30.0200 29.9000 30.1600 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1717 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5655 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met1  ;
    ANTENNAMAXAREACAR 14.2002 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 63.6354 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.27899 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.008 LAYER met2  ;
    ANTENNAGATEAREA 1.98 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7281 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.2151 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.27899 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 27.9800 29.9000 28.1200 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1973 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8415 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.431 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.98 LAYER met2  ;
    ANTENNAMAXAREACAR 11.8926 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.3247 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 26.9600 29.9000 27.1000 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1578 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5395 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 41.8083 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 203.901 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.846 LAYER met2  ;
    ANTENNAGATEAREA 1.737 LAYER met2  ;
    ANTENNAMAXAREACAR 45.8466 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 223.962 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 25.6000 29.9000 25.7400 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1985 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.878 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met1  ;
    ANTENNAMAXAREACAR 2.30626 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 8.26667 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.0540741 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8341 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8815 LAYER met2  ;
    ANTENNAGATEAREA 1.611 LAYER met2  ;
    ANTENNAMAXAREACAR 23.4154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.6078 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.840702 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAGATEAREA 1.611 LAYER met3  ;
    ANTENNAMAXAREACAR 23.835 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.1354 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.865532 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.44 LAYER met4  ;
    ANTENNAGATEAREA 1.737 LAYER met4  ;
    ANTENNAMAXAREACAR 54.4204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.291 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 23.9000 29.9000 24.0400 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3293 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.471 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 28.704 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 132.802 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.0988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.258 LAYER met2  ;
    ANTENNAGATEAREA 1.737 LAYER met2  ;
    ANTENNAMAXAREACAR 35.0936 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 164.614 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 22.5400 29.9000 22.6800 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.056 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.98 LAYER met1  ;
    ANTENNAMAXAREACAR 8.03318 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 20.2141 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.116768 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 20.8400 29.9000 20.9800 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9291 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.658 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.737 LAYER met2  ;
    ANTENNAMAXAREACAR 17.7147 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 43.6200 29.9000 43.7600 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1129 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.3085 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.611 LAYER met1  ;
    ANTENNAMAXAREACAR 4.99597 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 17.2495 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.243332 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3455 LAYER met2  ;
    ANTENNAGATEAREA 1.611 LAYER met2  ;
    ANTENNAMAXAREACAR 5.80497 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.1883 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.268161 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAGATEAREA 1.611 LAYER met3  ;
    ANTENNAMAXAREACAR 7.63799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.2541 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.29299 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.808 LAYER met4  ;
    ANTENNAGATEAREA 1.737 LAYER met4  ;
    ANTENNAMAXAREACAR 43.8936 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 41.9200 29.9000 42.0600 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2977 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 70.9937 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 333.365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 76.9063 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 368.603 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.912 LAYER met4  ;
    ANTENNAGATEAREA 1.737 LAYER met4  ;
    ANTENNAMAXAREACAR 82.783 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.216 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 40.5600 29.9000 40.7000 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.0768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.737 LAYER met4  ;
    ANTENNAMAXAREACAR 33.1585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.268 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.364707 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 38.8600 29.9000 39.0000 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6698 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.103 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.737 LAYER met1  ;
    ANTENNAMAXAREACAR 5.66206 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 20.5973 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 37.5000 29.9000 37.6400 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3005 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3205 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met1  ;
    ANTENNAMAXAREACAR 46.9631 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 104.002 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.548016 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met2  ;
    ANTENNAGATEAREA 1.737 LAYER met2  ;
    ANTENNAMAXAREACAR 48.6596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.416 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.548016 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 36.1400 29.9000 36.2800 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9277 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met1  ;
    ANTENNAMAXAREACAR 33.8444 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 156.956 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.0903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2805 LAYER met2  ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 74.2437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.728 LAYER met3  ;
    ANTENNAGATEAREA 1.737 LAYER met3  ;
    ANTENNAMAXAREACAR 75.0271 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 362.044 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 34.4400 29.9000 34.5800 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7963 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7655 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.3654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.473 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.989 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.0833 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.577778 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 29.3050 33.0800 29.9000 33.2200 ;
    END
  END W2END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 61.6400 29.9000 61.7800 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 59.9400 29.9000 60.0800 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 58.5800 29.9000 58.7200 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 57.2200 29.9000 57.3600 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 55.5200 29.9000 55.6600 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 54.1600 29.9000 54.3000 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 52.4600 29.9000 52.6000 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 51.1000 29.9000 51.2400 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 49.4000 29.9000 49.5400 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 48.0400 29.9000 48.1800 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 46.6800 29.9000 46.8200 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 29.3050 44.9800 29.9000 45.1200 ;
    END
  END W6END[0]
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.718 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 109.9200 0.5950 110.0600 ;
    END
  END A_I_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2505 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.7998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.736 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 105.8400 0.5950 105.9800 ;
    END
  END A_T_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.35 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.541 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met1  ;
    ANTENNAMAXAREACAR 2.72408 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 4.75065 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 101.7600 0.5950 101.9000 ;
    END
  END A_O_top
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.931 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.6744 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 341.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.304 LAYER met4  ;
    ANTENNAMAXAREACAR 29.1124 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.781 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0570313 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.3400 0.0000 15.4800 0.4850 ;
    END
  END UserCLK
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2133 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 98.0200 0.5950 98.1600 ;
    END
  END B_I_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.2137 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 93.9400 0.5950 94.0800 ;
    END
  END B_T_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2417 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0635 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.6984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.05 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.066 LAYER met2  ;
    ANTENNAMAXAREACAR 5.98991 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.4263 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 90.2000 0.5950 90.3400 ;
    END
  END B_O_top
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.45212 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.3892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 214.8400 0.8000 215.1400 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 9.9332 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.9279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 211.7900 0.8000 212.0900 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.16808 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.6364 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 208.7400 0.8000 209.0400 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.0638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2101 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 189.538 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.6900 0.8000 205.9900 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 33.5001 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 158.956 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.50915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 202.6400 0.8000 202.9400 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 15.6523 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 52.637 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.25109 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 199.5900 0.8000 199.8900 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.0768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 39.4601 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.452 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 196.5400 0.8000 196.8400 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.9258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 48.855 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.276 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 193.4900 0.8000 193.7900 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8205 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.1192 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 190.4400 0.8000 190.7400 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.87313 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.7104 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 187.3900 0.8000 187.6900 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.94101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.3717 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 184.3400 0.8000 184.6400 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 5.37791 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 25.0936 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 181.2900 0.8000 181.5900 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 19.4368 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 54.9597 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.25109 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 178.2400 0.8000 178.5400 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 12.4478 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.4767 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.367641 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 175.1900 0.8000 175.4900 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 30.5353 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.724 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.29546 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.1400 0.8000 172.4400 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.0248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 28.9172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.652 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 169.0900 0.8000 169.3900 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 6.74424 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.7279 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 166.0400 0.8000 166.3400 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.7188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.8651 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 292.329 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 162.9900 0.8000 163.2900 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 14.3573 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.5152 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 159.9400 0.8000 160.2400 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.90869 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.569 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 156.8900 0.8000 157.1900 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.53859 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.763 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 153.8400 0.8000 154.1400 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6636 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.0848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7547 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.358 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 150.7900 0.8000 151.0900 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 32.992 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.878 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.477221 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 147.7400 0.8000 148.0400 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.0918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met4  ;
    ANTENNAMAXAREACAR 35.1518 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.838 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 144.6900 0.8000 144.9900 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.9308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.9522 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.189 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 141.6400 0.8000 141.9400 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 2.15003 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 9.27677 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 138.5900 0.8000 138.8900 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.0296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.4676 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.864 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 135.5400 0.8000 135.8400 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 15.2752 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.5354 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 132.4900 0.8000 132.7900 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6526 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.9718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.5375 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.939 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 129.4400 0.8000 129.7400 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.467025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.5183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 48.3488 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 126.3900 0.8000 126.6900 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 21.3588 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.8169 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.25109 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 123.3400 0.8000 123.6400 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 19.1093 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.2287 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.50915 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 120.2900 0.8000 120.5900 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 214.8400 29.9000 215.1400 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 211.7900 29.9000 212.0900 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 208.7400 29.9000 209.0400 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.2956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 205.6900 29.9000 205.9900 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.472 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 202.6400 29.9000 202.9400 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 199.5900 29.9000 199.8900 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.224 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 196.5400 29.9000 196.8400 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 193.4900 29.9000 193.7900 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 190.4400 29.9000 190.7400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 187.3900 29.9000 187.6900 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7524 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 184.3400 29.9000 184.6400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.5798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.896 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 181.2900 29.9000 181.5900 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 178.2400 29.9000 178.5400 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 175.1900 29.9000 175.4900 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.8758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.808 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 172.1400 29.9000 172.4400 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 169.0900 29.9000 169.3900 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 166.0400 29.9000 166.3400 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.912 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 162.9900 29.9000 163.2900 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 159.9400 29.9000 160.2400 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 156.8900 29.9000 157.1900 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 153.8400 29.9000 154.1400 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.5546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.232 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 150.7900 29.9000 151.0900 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 147.7400 29.9000 148.0400 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4572 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 144.6900 29.9000 144.9900 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 141.6400 29.9000 141.9400 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 138.5900 29.9000 138.8900 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 135.5400 29.9000 135.8400 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.384 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 132.4900 29.9000 132.7900 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.608 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 129.4400 29.9000 129.7400 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 126.3900 29.9000 126.6900 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.136 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 123.3400 29.9000 123.6400 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9286 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.9458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.848 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 29.1000 120.2900 29.9000 120.5900 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.92 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.5428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 47.1134 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.276 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 26.8400 0.0000 26.9800 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.66828 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.365 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 0.0000 24.6800 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.87461 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.9919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 22.2400 0.0000 22.3800 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.167 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.871 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.4638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.0459 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.646 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 19.9400 0.0000 20.0800 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.1067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.426 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 38.596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 191.599 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 17.6400 0.0000 17.7800 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.3756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.374 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 331.331 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 13.0400 0.0000 13.1800 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.35542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.3461 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 10.7400 0.0000 10.8800 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2688 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.2411 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 8.4400 0.0000 8.5800 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2244 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.843 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.7786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8361 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.353 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 5.6800 0.0000 5.8200 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.06438 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.1805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 3.8400 0.0000 3.9800 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.2928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8238 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.3064 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 0.0000 27.9150 0.3300 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.7384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.574 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.7017 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.3407 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 0.0000 24.6950 0.3300 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.936 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.4664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.804 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 0.0000 21.9350 0.3300 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7584 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.718 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 5.98088 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 26.2923 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 0.0000 19.1750 0.3300 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.626 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.93253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.8061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 0.0000 16.4150 0.3300 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.3658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.8074 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.401 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 13.0250 0.0000 13.1950 0.3300 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.47 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.276 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 4.9697 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 23.6175 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.438 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.0435 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.4418 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 7.5050 0.0000 7.6750 0.3300 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.40345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.357 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.158 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 3.94451 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 16.1104 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 4.7450 0.0000 4.9150 0.3300 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.1987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.7045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1848 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.3258 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123707 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 12.2521 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.938 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.145265 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 15.8949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.4712 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.423899 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 1.9850 0.0000 2.1550 0.3300 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.7088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.584 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 26.3800 229.3550 26.5200 229.8400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.1888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 24.0800 229.3550 24.2200 229.8400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.894 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 248.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 21.3200 229.3550 21.4600 229.8400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5565 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.0200 229.3550 19.1600 229.8400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.5135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.2600 229.3550 16.4000 229.8400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.5000 229.3550 13.6400 229.8400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.2000 229.3550 11.3400 229.8400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.4400 229.3550 8.5800 229.8400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.6800 229.3550 5.8200 229.8400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.8197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.8725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.3800 229.3550 3.5200 229.8400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.3018 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.061 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.7336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 229.5100 27.9150 229.8400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.53645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.337 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.5284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.524 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.5250 229.5100 24.6950 229.8400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2486 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.469 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 229.5100 21.9350 229.8400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.38005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.153 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.595 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.472 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.0050 229.5100 19.1750 229.8400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8856 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6319 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.52 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 229.5100 16.4150 229.8400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.0250 229.5100 13.1950 229.8400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.242 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 229.5100 10.4350 229.8400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2304 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 7.5050 229.5100 7.6750 229.8400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.5932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.855 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 4.7450 229.5100 4.9150 229.8400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.7456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.584 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 1.9850 229.5100 2.1550 229.8400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 24.9100 5.4300 26.4100 224.0700 ;
        RECT 3.4900 5.4300 4.9900 224.0700 ;
      LAYER met3 ;
        RECT 3.4900 5.4300 26.4100 6.9300 ;
        RECT 3.4900 222.5700 26.4100 224.0700 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 27.4100 2.9300 28.9100 226.5700 ;
        RECT 0.9900 2.9300 2.4900 226.5700 ;
      LAYER met3 ;
        RECT 0.9900 2.9300 28.9100 4.4300 ;
        RECT 0.9900 225.0700 28.9100 226.5700 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 28.0850 229.3400 29.9000 229.8400 ;
      RECT 24.8650 229.3400 27.5750 229.8400 ;
      RECT 22.1050 229.3400 24.3550 229.8400 ;
      RECT 19.3450 229.3400 21.5950 229.8400 ;
      RECT 16.5850 229.3400 18.8350 229.8400 ;
      RECT 13.3650 229.3400 16.0750 229.8400 ;
      RECT 10.6050 229.3400 12.8550 229.8400 ;
      RECT 7.8450 229.3400 10.0950 229.8400 ;
      RECT 5.0850 229.3400 7.3350 229.8400 ;
      RECT 2.3250 229.3400 4.5750 229.8400 ;
      RECT 0.0000 229.3400 1.8150 229.8400 ;
      RECT 0.0000 0.5000 29.9000 229.3400 ;
      RECT 28.0850 0.0000 29.9000 0.5000 ;
      RECT 24.8650 0.0000 27.5750 0.5000 ;
      RECT 22.1050 0.0000 24.3550 0.5000 ;
      RECT 19.3450 0.0000 21.5950 0.5000 ;
      RECT 16.5850 0.0000 18.8350 0.5000 ;
      RECT 13.3650 0.0000 16.0750 0.5000 ;
      RECT 10.6050 0.0000 12.8550 0.5000 ;
      RECT 7.8450 0.0000 10.0950 0.5000 ;
      RECT 5.0850 0.0000 7.3350 0.5000 ;
      RECT 2.3250 0.0000 4.5750 0.5000 ;
      RECT 0.0000 0.0000 1.8150 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 110.2000 29.9000 229.8400 ;
      RECT 0.7350 109.8600 29.9000 110.2000 ;
      RECT 0.7350 109.7800 29.1650 109.8600 ;
      RECT 0.0000 109.4400 29.1650 109.7800 ;
      RECT 0.0000 108.5000 29.9000 109.4400 ;
      RECT 0.0000 108.0800 29.1650 108.5000 ;
      RECT 0.0000 107.1400 29.9000 108.0800 ;
      RECT 0.0000 106.7200 29.1650 107.1400 ;
      RECT 0.0000 106.1200 29.9000 106.7200 ;
      RECT 0.7350 105.7000 29.9000 106.1200 ;
      RECT 0.0000 105.4400 29.9000 105.7000 ;
      RECT 0.0000 105.0200 29.1650 105.4400 ;
      RECT 0.0000 104.0800 29.9000 105.0200 ;
      RECT 0.0000 103.6600 29.1650 104.0800 ;
      RECT 0.0000 102.3800 29.9000 103.6600 ;
      RECT 0.0000 102.0400 29.1650 102.3800 ;
      RECT 0.7350 101.9600 29.1650 102.0400 ;
      RECT 0.7350 101.6200 29.9000 101.9600 ;
      RECT 0.0000 101.0200 29.9000 101.6200 ;
      RECT 0.0000 100.6000 29.1650 101.0200 ;
      RECT 0.0000 99.3200 29.9000 100.6000 ;
      RECT 0.0000 98.9000 29.1650 99.3200 ;
      RECT 0.0000 98.3000 29.9000 98.9000 ;
      RECT 0.7350 97.9600 29.9000 98.3000 ;
      RECT 0.7350 97.8800 29.1650 97.9600 ;
      RECT 0.0000 97.5400 29.1650 97.8800 ;
      RECT 0.0000 96.6000 29.9000 97.5400 ;
      RECT 0.0000 96.1800 29.1650 96.6000 ;
      RECT 0.0000 94.9000 29.9000 96.1800 ;
      RECT 0.0000 94.4800 29.1650 94.9000 ;
      RECT 0.0000 94.2200 29.9000 94.4800 ;
      RECT 0.7350 93.8000 29.9000 94.2200 ;
      RECT 0.0000 93.5400 29.9000 93.8000 ;
      RECT 0.0000 93.1200 29.1650 93.5400 ;
      RECT 0.0000 91.8400 29.9000 93.1200 ;
      RECT 0.0000 91.4200 29.1650 91.8400 ;
      RECT 0.0000 90.4800 29.9000 91.4200 ;
      RECT 0.7350 90.0600 29.1650 90.4800 ;
      RECT 0.0000 88.7800 29.9000 90.0600 ;
      RECT 0.0000 88.3600 29.1650 88.7800 ;
      RECT 0.0000 87.4200 29.9000 88.3600 ;
      RECT 0.0000 87.0000 29.1650 87.4200 ;
      RECT 0.0000 86.0600 29.9000 87.0000 ;
      RECT 0.0000 85.6400 29.1650 86.0600 ;
      RECT 0.0000 84.3600 29.9000 85.6400 ;
      RECT 0.0000 83.9400 29.1650 84.3600 ;
      RECT 0.0000 83.0000 29.9000 83.9400 ;
      RECT 0.0000 82.5800 29.1650 83.0000 ;
      RECT 0.0000 81.3000 29.9000 82.5800 ;
      RECT 0.0000 80.8800 29.1650 81.3000 ;
      RECT 0.0000 79.9400 29.9000 80.8800 ;
      RECT 0.0000 79.5200 29.1650 79.9400 ;
      RECT 0.0000 78.2400 29.9000 79.5200 ;
      RECT 0.0000 77.8200 29.1650 78.2400 ;
      RECT 0.0000 76.8800 29.9000 77.8200 ;
      RECT 0.0000 76.4600 29.1650 76.8800 ;
      RECT 0.0000 75.5200 29.9000 76.4600 ;
      RECT 0.0000 75.1000 29.1650 75.5200 ;
      RECT 0.0000 73.8200 29.9000 75.1000 ;
      RECT 0.0000 73.4000 29.1650 73.8200 ;
      RECT 0.0000 72.4600 29.9000 73.4000 ;
      RECT 0.0000 72.0400 29.1650 72.4600 ;
      RECT 0.0000 70.7600 29.9000 72.0400 ;
      RECT 0.0000 70.3400 29.1650 70.7600 ;
      RECT 0.0000 69.4000 29.9000 70.3400 ;
      RECT 0.0000 68.9800 29.1650 69.4000 ;
      RECT 0.0000 67.7000 29.9000 68.9800 ;
      RECT 0.0000 67.2800 29.1650 67.7000 ;
      RECT 0.0000 66.3400 29.9000 67.2800 ;
      RECT 0.0000 65.9200 29.1650 66.3400 ;
      RECT 0.0000 64.9800 29.9000 65.9200 ;
      RECT 0.0000 64.5600 29.1650 64.9800 ;
      RECT 0.0000 63.2800 29.9000 64.5600 ;
      RECT 0.0000 62.8600 29.1650 63.2800 ;
      RECT 0.0000 61.9200 29.9000 62.8600 ;
      RECT 0.0000 61.5000 29.1650 61.9200 ;
      RECT 0.0000 60.2200 29.9000 61.5000 ;
      RECT 0.0000 59.8000 29.1650 60.2200 ;
      RECT 0.0000 58.8600 29.9000 59.8000 ;
      RECT 0.0000 58.4400 29.1650 58.8600 ;
      RECT 0.0000 57.5000 29.9000 58.4400 ;
      RECT 0.0000 57.0800 29.1650 57.5000 ;
      RECT 0.0000 55.8000 29.9000 57.0800 ;
      RECT 0.0000 55.3800 29.1650 55.8000 ;
      RECT 0.0000 54.4400 29.9000 55.3800 ;
      RECT 0.0000 54.0200 29.1650 54.4400 ;
      RECT 0.0000 52.7400 29.9000 54.0200 ;
      RECT 0.0000 52.3200 29.1650 52.7400 ;
      RECT 0.0000 51.3800 29.9000 52.3200 ;
      RECT 0.0000 50.9600 29.1650 51.3800 ;
      RECT 0.0000 49.6800 29.9000 50.9600 ;
      RECT 0.0000 49.2600 29.1650 49.6800 ;
      RECT 0.0000 48.3200 29.9000 49.2600 ;
      RECT 0.0000 47.9000 29.1650 48.3200 ;
      RECT 0.0000 46.9600 29.9000 47.9000 ;
      RECT 0.0000 46.5400 29.1650 46.9600 ;
      RECT 0.0000 45.2600 29.9000 46.5400 ;
      RECT 0.0000 44.8400 29.1650 45.2600 ;
      RECT 0.0000 43.9000 29.9000 44.8400 ;
      RECT 0.0000 43.4800 29.1650 43.9000 ;
      RECT 0.0000 42.2000 29.9000 43.4800 ;
      RECT 0.0000 41.7800 29.1650 42.2000 ;
      RECT 0.0000 40.8400 29.9000 41.7800 ;
      RECT 0.0000 40.4200 29.1650 40.8400 ;
      RECT 0.0000 39.1400 29.9000 40.4200 ;
      RECT 0.0000 38.7200 29.1650 39.1400 ;
      RECT 0.0000 37.7800 29.9000 38.7200 ;
      RECT 0.0000 37.3600 29.1650 37.7800 ;
      RECT 0.0000 36.4200 29.9000 37.3600 ;
      RECT 0.0000 36.0000 29.1650 36.4200 ;
      RECT 0.0000 34.7200 29.9000 36.0000 ;
      RECT 0.0000 34.3000 29.1650 34.7200 ;
      RECT 0.0000 33.3600 29.9000 34.3000 ;
      RECT 0.0000 32.9400 29.1650 33.3600 ;
      RECT 0.0000 31.6600 29.9000 32.9400 ;
      RECT 0.0000 31.2400 29.1650 31.6600 ;
      RECT 0.0000 30.3000 29.9000 31.2400 ;
      RECT 0.0000 29.8800 29.1650 30.3000 ;
      RECT 0.0000 28.2600 29.9000 29.8800 ;
      RECT 0.0000 27.8400 29.1650 28.2600 ;
      RECT 0.0000 27.2400 29.9000 27.8400 ;
      RECT 0.0000 26.8200 29.1650 27.2400 ;
      RECT 0.0000 25.8800 29.9000 26.8200 ;
      RECT 0.0000 25.4600 29.1650 25.8800 ;
      RECT 0.0000 24.1800 29.9000 25.4600 ;
      RECT 0.0000 23.7600 29.1650 24.1800 ;
      RECT 0.0000 22.8200 29.9000 23.7600 ;
      RECT 0.0000 22.4000 29.1650 22.8200 ;
      RECT 0.0000 21.1200 29.9000 22.4000 ;
      RECT 0.0000 20.7000 29.1650 21.1200 ;
      RECT 0.0000 19.7600 29.9000 20.7000 ;
      RECT 0.0000 19.3400 29.1650 19.7600 ;
      RECT 0.0000 18.0600 29.9000 19.3400 ;
      RECT 0.0000 17.6400 29.1650 18.0600 ;
      RECT 0.0000 16.7000 29.9000 17.6400 ;
      RECT 0.0000 16.2800 29.1650 16.7000 ;
      RECT 0.0000 15.3400 29.9000 16.2800 ;
      RECT 0.0000 14.9200 29.1650 15.3400 ;
      RECT 0.0000 0.0000 29.9000 14.9200 ;
    LAYER met2 ;
      RECT 26.6600 229.2150 29.9000 229.8400 ;
      RECT 24.3600 229.2150 26.2400 229.8400 ;
      RECT 21.6000 229.2150 23.9400 229.8400 ;
      RECT 19.3000 229.2150 21.1800 229.8400 ;
      RECT 16.5400 229.2150 18.8800 229.8400 ;
      RECT 13.7800 229.2150 16.1200 229.8400 ;
      RECT 11.4800 229.2150 13.3600 229.8400 ;
      RECT 8.7200 229.2150 11.0600 229.8400 ;
      RECT 5.9600 229.2150 8.3000 229.8400 ;
      RECT 3.6600 229.2150 5.5400 229.8400 ;
      RECT 0.0000 229.2150 3.2400 229.8400 ;
      RECT 0.0000 226.7100 29.9000 229.2150 ;
      RECT 2.6300 224.2100 27.2700 226.7100 ;
      RECT 26.5500 5.2900 27.2700 224.2100 ;
      RECT 5.1300 5.2900 24.7700 224.2100 ;
      RECT 2.6300 5.2900 3.3500 224.2100 ;
      RECT 29.0500 2.7900 29.9000 226.7100 ;
      RECT 2.6300 2.7900 27.2700 5.2900 ;
      RECT 0.0000 2.7900 0.8500 226.7100 ;
      RECT 0.0000 0.6250 29.9000 2.7900 ;
      RECT 27.1200 0.0000 29.9000 0.6250 ;
      RECT 24.8200 0.0000 26.7000 0.6250 ;
      RECT 22.5200 0.0000 24.4000 0.6250 ;
      RECT 20.2200 0.0000 22.1000 0.6250 ;
      RECT 17.9200 0.0000 19.8000 0.6250 ;
      RECT 15.6200 0.0000 17.5000 0.6250 ;
      RECT 13.3200 0.0000 15.2000 0.6250 ;
      RECT 11.0200 0.0000 12.9000 0.6250 ;
      RECT 8.7200 0.0000 10.6000 0.6250 ;
      RECT 5.9600 0.0000 8.3000 0.6250 ;
      RECT 4.1200 0.0000 5.5400 0.6250 ;
      RECT 0.0000 0.0000 3.7000 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 226.8700 29.9000 229.8400 ;
      RECT 29.2100 224.7700 29.9000 226.8700 ;
      RECT 0.0000 224.7700 0.6900 226.8700 ;
      RECT 0.0000 224.3700 29.9000 224.7700 ;
      RECT 26.7100 222.2700 29.9000 224.3700 ;
      RECT 0.0000 222.2700 3.1900 224.3700 ;
      RECT 0.0000 215.4400 29.9000 222.2700 ;
      RECT 1.1000 214.5400 28.8000 215.4400 ;
      RECT 0.0000 212.3900 29.9000 214.5400 ;
      RECT 1.1000 211.4900 28.8000 212.3900 ;
      RECT 0.0000 209.3400 29.9000 211.4900 ;
      RECT 1.1000 208.4400 28.8000 209.3400 ;
      RECT 0.0000 206.2900 29.9000 208.4400 ;
      RECT 1.1000 205.3900 28.8000 206.2900 ;
      RECT 0.0000 203.2400 29.9000 205.3900 ;
      RECT 1.1000 202.3400 28.8000 203.2400 ;
      RECT 0.0000 200.1900 29.9000 202.3400 ;
      RECT 1.1000 199.2900 28.8000 200.1900 ;
      RECT 0.0000 197.1400 29.9000 199.2900 ;
      RECT 1.1000 196.2400 28.8000 197.1400 ;
      RECT 0.0000 194.0900 29.9000 196.2400 ;
      RECT 1.1000 193.1900 28.8000 194.0900 ;
      RECT 0.0000 191.0400 29.9000 193.1900 ;
      RECT 1.1000 190.1400 28.8000 191.0400 ;
      RECT 0.0000 187.9900 29.9000 190.1400 ;
      RECT 1.1000 187.0900 28.8000 187.9900 ;
      RECT 0.0000 184.9400 29.9000 187.0900 ;
      RECT 1.1000 184.0400 28.8000 184.9400 ;
      RECT 0.0000 181.8900 29.9000 184.0400 ;
      RECT 1.1000 180.9900 28.8000 181.8900 ;
      RECT 0.0000 178.8400 29.9000 180.9900 ;
      RECT 1.1000 177.9400 28.8000 178.8400 ;
      RECT 0.0000 175.7900 29.9000 177.9400 ;
      RECT 1.1000 174.8900 28.8000 175.7900 ;
      RECT 0.0000 172.7400 29.9000 174.8900 ;
      RECT 1.1000 171.8400 28.8000 172.7400 ;
      RECT 0.0000 169.6900 29.9000 171.8400 ;
      RECT 1.1000 168.7900 28.8000 169.6900 ;
      RECT 0.0000 166.6400 29.9000 168.7900 ;
      RECT 1.1000 165.7400 28.8000 166.6400 ;
      RECT 0.0000 163.5900 29.9000 165.7400 ;
      RECT 1.1000 162.6900 28.8000 163.5900 ;
      RECT 0.0000 160.5400 29.9000 162.6900 ;
      RECT 1.1000 159.6400 28.8000 160.5400 ;
      RECT 0.0000 157.4900 29.9000 159.6400 ;
      RECT 1.1000 156.5900 28.8000 157.4900 ;
      RECT 0.0000 154.4400 29.9000 156.5900 ;
      RECT 1.1000 153.5400 28.8000 154.4400 ;
      RECT 0.0000 151.3900 29.9000 153.5400 ;
      RECT 1.1000 150.4900 28.8000 151.3900 ;
      RECT 0.0000 148.3400 29.9000 150.4900 ;
      RECT 1.1000 147.4400 28.8000 148.3400 ;
      RECT 0.0000 145.2900 29.9000 147.4400 ;
      RECT 1.1000 144.3900 28.8000 145.2900 ;
      RECT 0.0000 142.2400 29.9000 144.3900 ;
      RECT 1.1000 141.3400 28.8000 142.2400 ;
      RECT 0.0000 139.1900 29.9000 141.3400 ;
      RECT 1.1000 138.2900 28.8000 139.1900 ;
      RECT 0.0000 136.1400 29.9000 138.2900 ;
      RECT 1.1000 135.2400 28.8000 136.1400 ;
      RECT 0.0000 133.0900 29.9000 135.2400 ;
      RECT 1.1000 132.1900 28.8000 133.0900 ;
      RECT 0.0000 130.0400 29.9000 132.1900 ;
      RECT 1.1000 129.1400 28.8000 130.0400 ;
      RECT 0.0000 126.9900 29.9000 129.1400 ;
      RECT 1.1000 126.0900 28.8000 126.9900 ;
      RECT 0.0000 123.9400 29.9000 126.0900 ;
      RECT 1.1000 123.0400 28.8000 123.9400 ;
      RECT 0.0000 120.8900 29.9000 123.0400 ;
      RECT 1.1000 119.9900 28.8000 120.8900 ;
      RECT 0.0000 7.2300 29.9000 119.9900 ;
      RECT 26.7100 5.1300 29.9000 7.2300 ;
      RECT 0.0000 5.1300 3.1900 7.2300 ;
      RECT 0.0000 4.7300 29.9000 5.1300 ;
      RECT 29.2100 2.6300 29.9000 4.7300 ;
      RECT 0.0000 2.6300 0.6900 4.7300 ;
      RECT 0.0000 0.0000 29.9000 2.6300 ;
  END
END W_IO

END LIBRARY
